logic [23:0] sig_pr [0:12287] = {
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000000111111111111,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000001000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b111111111111000000000000,
24'b000000001100000000000101,
24'b000000000001000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000101,
24'b000000000001000000000000,
24'b000000001101000000000111,
24'b000000000000000000000001,
24'b000000001011000000000101,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000101,
24'b000000000001000000000000,
24'b000000001100000000000110,
24'b000000000000111111111111,
24'b000000001101000000000110,
24'b111111111111000000000001,
24'b000000001100000000000100,
24'b000000000001000000000000,
24'b000000001101000000000110,
24'b000000000000000000000001,
24'b000000001100000000000101,
24'b000000000000000000000001,
24'b000000001100000000000101,
24'b000000000001000000000001,
24'b000000001100000000000101,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b111111111111000000000000,
24'b000000001100000000000101,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b111111111111000000000000,
24'b000000001101000000000100,
24'b111111111111000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000001000000000001,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000001,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000001,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000001000000000000,
24'b000000001110000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000111111111111,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000000111111111111,
24'b000000001111000000000100,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000001000000000001,
24'b000000001110000000000100,
24'b000000000001000000000000,
24'b000000001111000000000100,
24'b000000000000000000000001,
24'b000000001110000000000100,
24'b111111111111000000000000,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001110000000000010,
24'b000000000000111111111111,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000010000000000000011,
24'b000000000000000000000000,
24'b000000001111000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000001000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000001000000000000,
24'b000000010000000000000011,
24'b000000000000000000000000,
24'b000000010001000000000010,
24'b000000000001000000000000,
24'b000000010001000000000011,
24'b000000000001000000000001,
24'b000000010000000000000011,
24'b000000000000000000000000,
24'b000000010000000000000011,
24'b111111111111000000000000,
24'b000000010001000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000000000000000000,
24'b000000010001000000000010,
24'b000000000000000000000000,
24'b000000010001000000000010,
24'b000000000000000000000000,
24'b000000010000000000000001,
24'b000000000000111111111111,
24'b000000010010000000000010,
24'b000000000000000000000001,
24'b000000010001000000000010,
24'b111111111111000000000000,
24'b000000010001000000000001,
24'b000000000000000000000000,
24'b000000010010000000000001,
24'b000000000000000000000000,
24'b000000010010000000000010,
24'b000000000000000000000000,
24'b000000010010000000000001,
24'b000000000000000000000001,
24'b000000010001000000000001,
24'b111111111111000000000000,
24'b000000010010000000000000,
24'b000000000000000000000001,
24'b000000010001000000000001,
24'b000000000000000000000000,
24'b000000010010000000000001,
24'b111111111111000000000000,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000001,
24'b000000000000000000000000,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000000,
24'b000000000000000000000001,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000000,
24'b000000000001000000000001,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000000,
24'b000000000001000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100111111111111,
24'b000000000001000000000000,
24'b000000010100000000000000,
24'b111111111111000000000000,
24'b000000010100111111111111,
24'b000000000000000000000000,
24'b000000010100111111111111,
24'b000000000001000000000000,
24'b000000010100000000000000,
24'b111111111111000000000000,
24'b000000010100111111111111,
24'b000000000001111111111111,
24'b000000010101000000000000,
24'b000000000000111111111111,
24'b000000010110111111111111,
24'b000000000000000000000000,
24'b000000010110111111111111,
24'b111111111111000000000000,
24'b000000010101111111111110,
24'b000000000001111111111111,
24'b000000010110111111111111,
24'b000000000000000000000000,
24'b000000010110111111111110,
24'b000000000000000000000000,
24'b000000010111111111111111,
24'b111111111111000000000000,
24'b000000010111111111111111,
24'b000000000000000000000000,
24'b000000010111111111111111,
24'b111111111111000000000000,
24'b000000010111111111111110,
24'b111111111111111111111111,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011001111111111110,
24'b000000000000000000000001,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011001111111111101,
24'b000000000000000000000000,
24'b000000011001111111111101,
24'b000000000000000000000000,
24'b000000011010111111111101,
24'b000000000000000000000000,
24'b000000011001111111111101,
24'b000000000001111111111111,
24'b000000011010111111111110,
24'b000000000000000000000000,
24'b000000011011111111111101,
24'b111111111111000000000000,
24'b000000011011111111111100,
24'b000000000000000000000001,
24'b000000011010111111111101,
24'b000000000000111111111111,
24'b000000011100111111111101,
24'b000000000000000000000000,
24'b000000011100111111111101,
24'b000000000000000000000000,
24'b000000011100111111111101,
24'b111111111111000000000000,
24'b000000011101111111111100,
24'b000000000000000000000000,
24'b000000011101111111111101,
24'b111111111111000000000000,
24'b000000011110111111111100,
24'b000000000000000000000000,
24'b000000011110111111111101,
24'b111111111111000000000000,
24'b000000011111111111111100,
24'b111111111111000000000000,
24'b000000011111111111111011,
24'b000000000000000000000000,
24'b000000100000111111111011,
24'b000000000000000000000001,
24'b000000100000111111111100,
24'b000000000000000000000000,
24'b000000100001111111111011,
24'b000000000000000000000000,
24'b000000100001111111111011,
24'b000000000000000000000000,
24'b000000100010111111111011,
24'b000000000000000000000001,
24'b000000100010111111111011,
24'b000000000000000000000000,
24'b000000100011111111111010,
24'b000000000000000000000000,
24'b000000100100111111111011,
24'b111111111111000000000000,
24'b000000100101111111111010,
24'b111111111111000000000000,
24'b000000100110111111111001,
24'b000000000000000000000001,
24'b000000100110111111111010,
24'b000000000000000000000000,
24'b000000100111111111111010,
24'b000000000000000000000000,
24'b000000101001111111111010,
24'b000000000000000000000001,
24'b000000101001111111111010,
24'b111111111111000000000000,
24'b000000101010111111111001,
24'b111111111111000000000000,
24'b000000101010111111111000,
24'b000000000000111111111111,
24'b000000101100111111111001,
24'b111111111111111111111111,
24'b000000101110111111111000,
24'b000000000000000000000000,
24'b000000101111111111111000,
24'b111111111111000000000000,
24'b000000110001111111111000,
24'b000000000000000000000001,
24'b000000110001111111110111,
24'b000000000000000000000000,
24'b000000110011111111110111,
24'b000000000000000000000000,
24'b000000110101111111110110,
24'b000000000000000000000000,
24'b000000110111111111110110,
24'b000000000000000000000001,
24'b000000111000111111110110,
24'b000000000000000000000000,
24'b000000111011111111110110,
24'b000000000000000000000001,
24'b000000111101111111110101,
24'b000000000000000000000000,
24'b000000111110111111110101,
24'b000000000000111111111111,
24'b000001000011111111110100,
24'b000000000000000000000000,
24'b000001000110111111110100,
24'b000000000000000000000000,
24'b000001001001111111110011,
24'b000000000000000000000000,
24'b000001001100111111110010,
24'b000000000000000000000000,
24'b000001010001111111110000,
24'b000000000001000000000000,
24'b000001010101111111101111,
24'b000000000000111111111111,
24'b000001011011111111101110,
24'b111111111111000000000000,
24'b000001100001111111101010,
24'b000000000000000000000000,
24'b000001101001111111100111,
24'b111111111111000000000000,
24'b000001110000111111100010,
24'b000000000000000000000000,
24'b000001111010111111011011,
24'b000000000001000000000001,
24'b000010000100111111010001,
24'b000000000000000000000000,
24'b000010010000111111000000,
24'b000000000000000000000000,
24'b000010011100111110100000,
24'b000000000000000000000000,
24'b000010011010111101010110,
24'b000000000000000000000000,
24'b111111010111110111111011,
24'b001011010110110100101010,
24'b010100001011000010010110,
24'b001011010110001011010110,
24'b000110111001010000001110,
24'b110100101010001011010110,
24'b000001000111111000000011,
24'b001011010110001011010110,
24'b110101000100001110010001,
24'b110100101001110100101001,
24'b010000000010110111100000,
24'b001011010101001011010101,
24'b000100101001001110011010,
24'b110100101001001011010110,
24'b000000110111111000010101,
24'b001011010101001011010101,
24'b111101111000010000100110,
24'b110100101010001011010110,
24'b111010000010000010100110,
24'b110100101010001011010110,
24'b101110011101110101000000,
24'b001011010101110100101010,
24'b001001000001001111000111,
24'b110100101010001011010110,
24'b111011110101000010111011,
24'b110100101001001011010111,
24'b101110010011111110000010,
24'b110100101010110100101010,
24'b000111101111111000110001,
24'b110100101010001011010110,
24'b111001010001101010110000,
24'b001011010110001011010110,
24'b101001010001111010100110,
24'b001011010110110100101010,
24'b110111101101000010110011,
24'b001011010110110100101001,
24'b111101100110010010100111,
24'b110100101011110100101010,
24'b000011011000000100100010,
24'b110100101001110100101010,
24'b010001011101111111000111,
24'b110100101010001011010101,
24'b000000101100111010000011,
24'b110100101010001011010101,
24'b110000010011101101100100,
24'b001011010101110100101010,
24'b000000000010000111001010,
24'b110100101011110100101010,
24'b001111010010111000101011,
24'b110100101010001011010111,
24'b111000001110101000100010,
24'b001011010110110100101010,
24'b010000100001110110110010,
24'b001011010110001011010110,
24'b000011100010111100011000,
24'b001011010110001011010111,
24'b111110001100000001101001,
24'b001011010110001011010110,
24'b111000100110001110011101,
24'b110100101001001011010110,
24'b101010010001110101110010,
24'b001011010110110100101010,
24'b111001110011001011101001,
24'b110100101001110100101011,
24'b000001100000110100100001,
24'b001011010110110100101010,
24'b010000100000001010111111,
24'b110100101010001011010110,
24'b000000100001110100001100,
24'b001011010110001011010101,
24'b110001100011001010111010,
24'b110100101010110100101010,
24'b001001011011110100100001,
24'b001011010110001011010110,
24'b110011010000001100010100,
24'b110100101010110100101010,
24'b001010011001111101100011,
24'b110100101010001011010110,
24'b110100010111101110101001,
24'b001011010110110100101010,
24'b001100101011000101111101,
24'b110100101011001011010110,
24'b111111000101101110001010,
24'b001011010110001011010110,
24'b110111111011111100100000,
24'b001011010110001011010111,
24'b101000101011001010011110,
24'b110100101010110100101010,
24'b110111001010110000111111,
24'b001011010110110100101010,
24'b111100111001111110110011,
24'b001011010111110100101010,
24'b000010011010001100110101,
24'b110100101010110100101001,
24'b010000001010110100010100,
24'b001011010110001011010111,
24'b111110110100001001110110,
24'b110100101010001011010110,
24'b101101100011110001100001,
24'b001011010110110100101010,
24'b111011011011000000000001,
24'b001011010110110100101010,
24'b000001101101001111011000,
24'b110100101010110100101010,
24'b001110011100111110111111,
24'b110100101011001011010101,
24'b110100101111101111010001,
24'b001011010110110100101001,
24'b000010110111000101110111,
24'b110100101010110100101001,
24'b010010001001101101001001,
24'b001011010111001011010101,
24'b000001111010111001100111,
24'b001011010110001011010110,
24'b110010011111111110001101,
24'b001011010111110100101010,
24'b001001101011000010101000,
24'b001011010110001011011000,
24'b110001111110001110011001,
24'b110100101010110100101010,
24'b000000110101110011101110,
24'b001011010110110100101010,
24'b010000010110000000000001,
24'b001011010110001011010110,
24'b111111110110000110001100,
24'b001011010111001011010110,
24'b101111001010010100011100,
24'b110100101010110100101010,
24'b111101101110000100100111,
24'b110100101010110100101010,
24'b000101000100111100011010,
24'b110100101001110100101010,
24'b010100001100101100100011,
24'b001011010110001011010110,
24'b000101011010111010101010,
24'b001011010111001011010111,
24'b111111001010000000001011,
24'b001011010111001011010110,
24'b111000110100000101101000,
24'b001011010110001011010111,
24'b101001101001010011011101,
24'b110100101010110100101010,
24'b110111111011000010100110,
24'b110100101010110100101011,
24'b111101000011110010110010,
24'b001011010111110100101010,
24'b000000111100001001101001,
24'b110100101010110100101010,
24'b000101011111110001100011,
24'b001011010110110100101010,
24'b010001110110111111101110,
24'b001011010101001011010110,
24'b111000101111001101101000,
24'b110100101010110100101001,
24'b001101111101110100001111,
24'b001011010110001011010110,
24'b110101010000000010011000,
24'b001011010110110100101001,
24'b000010101100010001100000,
24'b110100101010110100101011,
24'b001001110101000000110001,
24'b110100101010110100101010,
24'b011001001110110000000011,
24'b001011010110001011010110,
24'b001011000110111111001011,
24'b001011010110001011010110,
24'b000110001100001101010011,
24'b110100101001001011010110,
24'b000010110001110011110111,
24'b001011010101001011010110,
24'b111111011111000001101010,
24'b001011010101001011010111,
24'b111011000011001111100001,
24'b110100101010001011010111,
24'b101110000000110110010100,
24'b001011010101110100101010,
24'b111111110110000100110110,
24'b001011010110110100101010,
24'b010001101011010100110011,
24'b110100101010001011010110,
24'b000100101000000110000101,
24'b110100101010001011010110,
24'b000000001101111111001101,
24'b110100101010001011010101,
24'b111100111101110001111011,
24'b001011010110001011010101,
24'b111001100100001011001001,
24'b110100101011001011010110,
24'b110100110000111100011110,
24'b110100101001001011010110,
24'b100110111001101100010111,
24'b001011010110110100101010,
24'b110111010000111011000001,
24'b001011010110110100101011,
24'b000101110110000010000101,
24'b001011010110001011010110,
24'b101100010010010000011001,
24'b110100101011110100101010,
24'b111000111000111111011101,
24'b110100101010110100101010,
24'b111110100000101110100110,
24'b001011010110110100101001,
24'b001010100101111101100101,
24'b001011010101001011010110,
24'b101111101100001011011100,
24'b110100101010110100101010,
24'b111011001110110001100001,
24'b001011010110110100101010,
24'b111111001000111110000001,
24'b001011010110110100101010,
24'b000010010111000011111001,
24'b001011010101110100101010,
24'b000110100001010000101011,
24'b110100101010110100101001,
24'b010010101101110111110011,
24'b001011010110001011010110,
24'b111001100111001101011010,
24'b110100101001110100101010,
24'b001111001100110101111101,
24'b001011010101001011010110,
24'b110111111001001011111011,
24'b110100101010110100101010,
24'b001110010001110100011110,
24'b001011010110001011010110,
24'b110111100110001010000001,
24'b110100101010110100101010,
24'b001111000101110001000011,
24'b001011010110001011010110,
24'b111111110010111101100100,
24'b001011010110001011010111,
24'b101111011111000010100000,
24'b001011010110110100101010,
24'b111110001100000111101000,
24'b001011010111110100101010,
24'b000101100011010101010010,
24'b110100101010110100101010,
24'b010100100011000100001010,
24'b110100101010001011010110,
24'b000101011000110011100011,
24'b001011010110001011010101,
24'b111101111000000011010011,
24'b001011010110001011010111,
24'b101110111101010011011010,
24'b110100101010110100101010,
24'b111110111101000100010110,
24'b110100101010110100101001,
24'b001101110011111100100000,
24'b110100101010001011010110,
24'b110101000110101100110011,
24'b001011010110110100101010,
24'b000011111111111010110100,
24'b001011010110110100101010,
24'b010100001010111111111001,
24'b001011010110001011010110,
24'b000101100110000011111000,
24'b001011010110001011010101,
24'b111110110010001000110000,
24'b001011010110001011010111,
24'b110001010110010110001111,
24'b110100101010110100101010,
24'b001001101101000100111100,
24'b110100101001001011010110,
24'b110011101010110011110111,
24'b001011010110110100101010,
24'b001010101000000010001110,
24'b001011010110001011010110,
24'b110100000011001001011100,
24'b001011010110110100101010,
24'b001010101111011000010110,
24'b110100101010001011010110,
24'b110011111010001000101001,
24'b110100101010110100101010,
24'b001010001110111010100001,
24'b001011010110001011010110,
24'b110010010111010100100100,
24'b110100101010110100101010,
24'b000001001110001000101101,
24'b110100101010110100101010,
24'b010000110100000100110001,
24'b110100101010001011010110,
24'b000000011111000001111000,
24'b110100101010001011010111,
24'b110000001001111111000000,
24'b110100101011110100101010,
24'b111111110001111011000110,
24'b110100101010110100101001,
24'b001110101110101111010010,
24'b001011010110001011010101,
24'b110111001001001001011100,
24'b110100101010110100101010,
24'b001110011010111011011011,
24'b110100101010001011010110,
24'b111111000101101011110111,
24'b001011010110001011010110,
24'b101110111100111010111011,
24'b001011010111110100101011,
24'b111110010111000010010001,
24'b001011010110110100101010,
24'b001100101101010000010011,
24'b110100101001001011010110,
24'b110011011010111000110101,
24'b001011010110110100101010,
24'b000001010001010000111001,
24'b110100101010110100101011,
24'b001111000110000011100111,
24'b110100101010001011010111,
24'b110101101101111101010111,
24'b110100101011110100101010,
24'b000011110011110000100001,
24'b001011010101110100101001,
24'b010010010100001010000010,
24'b110100101010001011010101,
24'b111010110010111011101010,
24'b110100101001110100101011,
24'b010010100011101011110111,
24'b001011010110001011010110,
24'b000100110101111010110111,
24'b001011010110001011010110,
24'b111101110101000010011010,
24'b001011010110001011010110,
24'b101111001100010001100010,
24'b110100101011110100101010,
24'b111111010101000010011111,
24'b110100101010110100101010,
24'b001110001100111011001010,
24'b110100101010001011010110,
24'b110101011101101101000100,
24'b001011010110110100101010,
24'b000100001100000100010010,
24'b110100101011110100101010,
24'b010011111001101011110101,
24'b001011010111001011010101,
24'b000011111000111000010011,
24'b001011010110001011010110,
24'b110100000110111100100100,
24'b001011010110110100101010,
24'b000100101001111111110110,
24'b001011010110110100101010,
24'b010101101011000011101101,
24'b001011010110001011010111,
24'b000111111011001111000101,
24'b110100101010001011010110,
24'b000010100110110011111011,
24'b001011010110001011010110,
24'b111101010011111111011101,
24'b001011010111001011010110,
24'b101111101101000011101111,
24'b001011010110110100101010,
24'b000000111111001000001111,
24'b001011010110110100101010,
24'b010010000000010100100101,
24'b110100101011001011010101,
24'b000011000001111011100111,
24'b001011010110001011010110,
24'b110100110101010001010001,
24'b110100101010110100101011,
24'b001101011101111010000100,
24'b001011010110001011010101,
24'b111000011000010000100001,
24'b110100101010110100101010,
24'b010001100110111001110101,
24'b001011010101001011010110,
24'b000101001010010000110000,
24'b110100101010001011010101,
24'b111111110001111010110000,
24'b001011010110001011010110,
24'b110011111010010011010010,
24'b110100101010110100101011,
24'b001110111100000110001100,
24'b110100101010001011010110,
24'b000011100100000000000010,
24'b110100101010001011010110,
24'b111111101101110011000101,
24'b001011010110001011010110,
24'b111100011100001011111110,
24'b110100101010001011010101,
24'b111000000010110110101001,
24'b001011010111001011010110,
24'b101010110011001111010000,
24'b110100101010110100101010,
24'b111100000100000001010010,
24'b110100101010110100101010,
24'b001100001100110011011100,
24'b001011010110001011010110,
24'b110101101101001100111010,
24'b110100101010110100101010,
24'b001110010101111110111101,
24'b110100101010001011010111,
24'b000001010110110000101011,
24'b001011010110001011010110,
24'b111011010010001000101011,
24'b110100101010001011010110,
24'b101110010110110010001110,
24'b001011010110110100101010,
24'b000111000100001000011100,
24'b110100101011001011010110,
24'b110001010011101111111111,
24'b001011010111110100101010,
24'b001000100000111100111011,
24'b001011010110001011010110,
24'b110010000111000010001011,
24'b001011010110110100101001,
24'b001000110101000111100001,
24'b001011010110001011010110,
24'b110001011011010100110010,
24'b110100101010110100101010,
24'b000000110101111101000101,
24'b001011010110110100101010,
24'b010001010100010101001101,
24'b110100101010001011010110,
24'b000010111010001000011110,
24'b110100101010001011010110,
24'b111100000010000011111101,
24'b110100101011001011010110,
24'b101101110111000000100011,
24'b110100101010110100101010,
24'b111111000001111101000010,
24'b110100101010110100101001,
24'b010000010100111000000101,
24'b110100101010001011010111,
24'b000010100111101001111110,
24'b001011010110001011010110,
24'b111101001101111001011010,
24'b001011010110001011010111,
24'b110111101101000000100111,
24'b001011010110001011010111,
24'b101001101100001110000010,
24'b110100101011110100101010,
24'b111010010001110100110110,
24'b001011010110110100101010,
24'b001001100110000011011010,
24'b001011010110001011010101,
24'b110001111111010011001011,
24'b110100101001110100101010,
24'b001000010011000011011110,
24'b110100101010001011010110,
24'b110001010000110100111010,
24'b001011010110110100101001,
24'b000111011000001101111111,
24'b110100101010001011010111,
24'b101111001101111111110000,
24'b110100101010110100101010,
24'b111101011111110001001110,
24'b001011010110110100101010,
24'b001011100100001000111000,
24'b110100101010001011010110,
24'b110010010111110001011100,
24'b001011010110110100101010,
24'b000000101111000000001011,
24'b001011010110110100101010,
24'b010000001010001110101011,
24'b110100101001001011010110,
24'b111111111110110101111011,
24'b001011010110001011010101,
24'b110000100011000100111100,
24'b001011010111110100101010,
24'b000111100101010101011100,
24'b110100101001001011010110,
24'b101111011110000111100000,
24'b110100101001110100101001,
24'b111101000000000010010100,
24'b110100101010110100101010,
24'b000011110101111110000110,
24'b110100101010110100101010,
24'b010010011000111000101111,
24'b110100101011001011010110,
24'b000010001000101010010110,
24'b001011010110001011010110,
24'b110011000001111001011001,
24'b001011010110110100101010,
24'b001010111011111111100111,
24'b001011010110001011010110,
24'b110101000101000101101011,
24'b001011010101110100101010,
24'b001101011101010100000110,
24'b110100101010001011010110,
24'b111111111011000011111010,
24'b110100101001001011010110,
24'b111000110101110100111010,
24'b001011010110001011010110,
24'b101001110001001100111101,
24'b110100101010110100101010,
24'b111000101001110111001111,
24'b001011010111110100101010,
24'b111111100001001111101011,
24'b110100101001110100101010,
24'b001100110101000001101000,
24'b110100101010001011010110,
24'b110100001100110011111011,
24'b001011010110110100101010,
24'b001001101100001101110001,
24'b110100101001001011010101,
24'b110001010011000000111110,
24'b110100101010110100101011,
24'b111111100011111010100011,
24'b110100101001110100101100,
24'b001101111001101100010101,
24'b001011010111001011010110,
24'b110101111110111101000100,
24'b001011010110110100101010,
24'b001100111100001101010100,
24'b110100101010001011010101,
24'b111101010100111101001001,
24'b110100101010001011010110,
24'b101100101010101100011111,
24'b001011010110110100101010,
24'b111010111001111010110001,
24'b001011010111110100101011,
24'b000001011011000001010111,
24'b001011010111110100101010,
24'b001110100011001110011110,
24'b110100101010001011010110,
24'b110101111001110101100111,
24'b001011010111110100101011,
24'b001011100010001010110001,
24'b110100101010001011010110,
24'b110100000011110001101100,
24'b001011010111110100101010,
24'b001001101111111110001111,
24'b001011010110001011010110,
24'b110001000101000011001100,
24'b001011010111110100101010,
24'b111110010011001000010010,
24'b001011010110110100101010,
24'b000100111110010101010001,
24'b110100101011110100101011,
24'b010011100001111101001100,
24'b001011010110001011010110,
24'b000011111100010100101010,
24'b110100101010001011010110,
24'b111011111011000110010000,
24'b110100101010001011010110,
24'b101100010010111000100000,
24'b001011010110110100101010,
24'b111010101110010010100110,
24'b110100101010110100101010,
24'b000001001001000110100101,
24'b110100101011110100101010,
24'b001101110001000010010000,
24'b110100101010001011010101,
24'b110011100110111110100001,
24'b110100101010110100101010,
24'b000000001110111001100100,
24'b110100101010110100101010,
24'b000110100110101011100100,
24'b001011010111110100101010,
24'b010100110111111011001101,
24'b001011010111001011010111,
24'b000100011011000010110000,
24'b001011010101001011010101,
24'b110101010111010000101110,
24'b110100101010110100101010,
24'b001101111010111000111100,
24'b001011010101001011010110,
24'b111111000000001111100111,
24'b110100101010001011010110,
24'b101111000010111001100100,
24'b001011010111110100101010,
24'b111110100101010001111101,
24'b110100101010110100101010,
24'b001100111111000100000011,
24'b110100101010001011010110,
24'b110011110001110110100001,
24'b001011010110110100101010,
24'b000001110000010000100001,
24'b110100101010110100101010,
24'b001111110011000011011011,
24'b110100101010001011010110,
24'b110110110000110110100100,
24'b001011010110110100101010,
24'b000101011111010001011110,
24'b110100101010110100101001,
24'b010101101110000110010010,
24'b110100101011001011010110,
24'b000111011101000011000000,
24'b110100101010001011010110,
24'b000001101110000000110110,
24'b110100101001001011010110,
24'b111100000101111111000010,
24'b110100101010001011010101,
24'b101110001000111101010011,
24'b110100101010110100101010,
24'b111111000010111011011000,
24'b110100101010110100101011,
24'b001111100010111000111110,
24'b110100101010001011010110,
24'b111111111101110101001100,
24'b110100101010001011010111,
24'b110000110110101001000101,
24'b001011010110110100101010,
24'b001000000101000001111000,
24'b110100101010001011010110,
24'b110000000101101011000100,
24'b001011010110110100101001,
24'b111101100100111010001101,
24'b001011010110110100101010,
24'b000100000111001001000001,
24'b110100101001110100101010,
24'b010001100011110000111101,
24'b001011010111001011010110,
24'b111001011001000110101110,
24'b110100101010110100101010,
24'b001111111011101110001101,
24'b001011010110001011010110,
24'b111001110111111011011111,
24'b001011010110110100101010,
24'b010010100111000010001001,
24'b001011010110001011010110,
24'b000110001010010000011000,
24'b110100101010001011010111,
24'b000001101111111111100010,
24'b110100101010001011010110,
24'b111110010101101110111100,
24'b001011010111001011010101,
24'b111010110001111110010110,
24'b001011010110001011010110,
24'b110101101011001101000001,
24'b110100101010001011010110,
24'b100111010100110100111010,
24'b001011010110110100101010,
24'b110110001111001010110001,
24'b110100101010110100101010,
24'b111100001111110010101101,
24'b001011010110110100101010,
24'b000001111000000001011111,
24'b001011010111110100101010,
24'b001111101010010001000101,
24'b110100101010001011010110,
24'b111110010101000000110011,
24'b110100101010001011010110,
24'b101100111110110000100111,
24'b001011010110110100101010,
24'b111010101010000000011010,
24'b001011010110110100101100,
24'b000000100100001111101001,
24'b110100101010110100101001,
24'b001100110000111000100010,
24'b001011010110001011010110,
24'b110001111011010000101000,
24'b110100101010110100101011,
24'b111101011100000011001101,
24'b110100101010110100101010,
24'b000001010101111100100010,
24'b110100101010110100101010,
24'b000100011000101110010101,
24'b001011010110110100101010,
24'b000111101010111111010000,
24'b001011010110110100101010,
24'b001100011011010000000001,
24'b110100101001110100101001,
24'b011010000101000001000010,
24'b110100101010001011010110,
24'b000110110100110101101111,
24'b000000000000000000000000,
24'b010000001111110110111100,
24'b001011010110001011010100,
24'b001000001011001010011101,
24'b110100101010001011010101,
24'b000100011110110010101100,
24'b001011010110001011010110,
24'b000001001110000001111011,
24'b001011010101001011010110,
24'b111101001000010010001000,
24'b110100101010001011010110,
24'b110001001010000010111000,
24'b110100101001110100101010,
24'b001010101100110100110101,
24'b001011010110001011010111,
24'b110110000000001110110000,
24'b110100101010110100101010,
24'b001111011110000010011100,
24'b110100101010001011010110,
24'b000011010101111101011111,
24'b110100101011001011010110,
24'b111110110101111000001001,
24'b110100101010001011010110,
24'b111010011000101010000011,
24'b001011010110001011010110,
24'b101110011011111001110101,
24'b001011010110110100101011,
24'b001000110011000001111000,
24'b001011010111001011010110,
24'b111100000010010001100100,
24'b110100101001001011010101,
24'b110101001111000011001011,
24'b110100101010001011010101,
24'b100110000010111101010111,
24'b110100101010110100101010,
24'b110100001100110111100000,
24'b110100101010110100101010,
24'b111001000110101001000101,
24'b001011010111110100101001,
24'b111100011011111001000101,
24'b001011010110110100101001,
24'b111111011100000111011011,
24'b110100101011110100101010,
24'b000011010000101101100111,
24'b001011010110110100101010,
24'b001110101000111001101101,
24'b001011010110001011010110,
24'b110011100010111101111111,
24'b001011010110110100101001,
24'b111111001010000001010010,
24'b001011010110110100101001,
24'b000011100100000100110011,
24'b001011010110110100101010,
24'b001000001110001001110100,
24'b001011010110110100101010,
24'b010100110100011000000011,
24'b110100101001001011010101,
24'b111100011000001000110001,
24'b110100101001110100101011,
24'b010011010111000001101110,
24'b110100101010001011010101,
24'b000100010110110100011101,
24'b001011010110001011010110,
24'b110101100010001101010011,
24'b110100101010110100101010,
24'b001101010111111000010010,
24'b001011010110001011010101,
24'b110111000011010001101001,
24'b110100101001110100101010,
24'b001101110000000101100111,
24'b110100101010001011010110,
24'b110110011010000001100110,
24'b110100101011110100101010,
24'b000110000010111110101001,
24'b110100101010110100101011,
24'b010110111011111011100011,
24'b110100101011001011010110,
24'b001001011011110111001100,
24'b110100101010001011010101,
24'b000100110101101001111101,
24'b001011010111001011010110,
24'b000001100011111011011000,
24'b001011010110001011010110,
24'b111110010011001100010001,
24'b110100101010001011010110,
24'b111001110101111100110111,
24'b110100101010001011010110,
24'b101100100101101101011000,
24'b001011010110110100101010,
24'b111110000010111110000100,
24'b001011010110110100101011,
24'b001111000100001111000101,
24'b110100101010001011010110,
24'b000000000100000001001100,
24'b110100101010001011010110,
24'b110001111000111011100011,
24'b110100101010110100101010,
24'b001011000100110101101110,
24'b110100101011001011010101,
24'b111100101011100111001100,
24'b001011010110001011010110,
24'b101101001100110110011000,
24'b001011010111110100101011,
24'b111101001111111101101011,
24'b001011010110110100101011,
24'b001100011010001100000001,
24'b110100101011001011010110,
24'b110100111100111010111010,
24'b110100101010110100101010,
24'b001100001011101001100000,
24'b001011010110001011010110,
24'b111100101000110110110110,
24'b001011010110001011010101,
24'b101011111011111011100000,
24'b001011010110110100101010,
24'b111001101100111111001010,
24'b001011010110110100101010,
24'b111110101011000011101101,
24'b001011010110110100101001,
24'b000010101000010000110100,
24'b110100101010110100101010,
24'b000111010111111110111111,
24'b110100101011110100101011,
24'b010100000011101101001011,
24'b001011010110001011010110,
24'b111011100010111010001111,
24'b001011010111110100101010,
24'b010001110110111110110000,
24'b001011010110001011010110,
24'b111011101001000010010001,
24'b001011010110110100101011,
24'b010100001101000110101000,
24'b001011010111001011010110,
24'b000111010110010010111101,
24'b110100101010001011010110,
24'b000001101000111010000001,
24'b001011010110001011010111,
24'b110101100100001111110010,
24'b110100101010110100101010,
24'b010000100000111000101100,
24'b001011010111001011010110,
24'b000101000101001111011001,
24'b110100101010001011010110,
24'b000001010010111001001000,
24'b001011010110001011010101,
24'b111110010000010001010011,
24'b110100101001001011010111,
24'b111010011000000011001010,
24'b110100101001001011010110,
24'b101110110010110101011101,
24'b001011010110110100101010,
24'b001001010100001111011111,
24'b110100101010001011010110,
24'b111100000111000011001111,
24'b110100101010001011010111,
24'b101110100101111110010100,
24'b110100101011110100101010,
24'b000111111111111001000001,
24'b110100101010001011010110,
24'b111001011111101010111100,
24'b001011010110001011010110,
24'b101001011111111010110001,
24'b001011010110110100101001,
24'b110111111011000010111011,
24'b001011010101110100101001,
24'b111101110100010010101101,
24'b110100101010110100101011,
24'b000011100100000100100101,
24'b110100101010110100101010,
24'b010001101010111111001010,
24'b110100101010001011010110,
24'b000000110111111010000101,
24'b110100101010001011010110,
24'b110000011101101101100100,
24'b001011010110110100101010,
24'b000000001100000111001010,
24'b110100101011110100101010,
24'b001111011010111000101001,
24'b110100101010001011010101,
24'b111000011000101000100001,
24'b001011010110110100101011,
24'b010000101000110110101111,
24'b001011010110001011010101,
24'b000011101010111100010100,
24'b001011010110001011010110,
24'b111110010101000001100100,
24'b001011010110001011010110,
24'b111000101110001110011000,
24'b110100101010001011010110,
24'b101010011000110101101101,
24'b001011010110110100101001,
24'b111001111010001011100011,
24'b110100101010110100101010,
24'b000001100111110100011100,
24'b001011010110110100101001,
24'b010000101000001010111000,
24'b110100101010001011010110,
24'b000000101000110100000101,
24'b001011010110001011010101,
24'b110001101011001010110010,
24'b110100101010110100101010,
24'b001001100001110100011001,
24'b001011010110001011010101,
24'b110011010111001100001100,
24'b110100101010110100101010,
24'b001010011111111101011010,
24'b110100101010001011010101,
24'b110100011111101110100000,
24'b001011010110110100101011,
24'b001100110001000101110100,
24'b110100101011001011010110,
24'b111111001100101110000001,
24'b001011010110001011010110,
24'b111000000000111100010111,
24'b001011010110001011010110,
24'b101000110001001010010100,
24'b110100101001110100101010,
24'b110111010000110000110101,
24'b001011010110110100101010,
24'b111100111111111110101001,
24'b001011010110110100101011,
24'b000010011111001100101010,
24'b110100101010110100101010,
24'b010000001110110100001001,
24'b001011010110001011010110,
24'b111110111010001001101011,
24'b110100101001001011010110,
24'b101101101000110001010101,
24'b001011010111110100101010,
24'b111011100000111111110111,
24'b001011010110110100101010,
24'b000001110001001111001101,
24'b110100101010110100101010,
24'b001110100010111110110100,
24'b110100101010001011010110,
24'b110100110101101111000100,
24'b001011010110110100101011,
24'b000010111011000101101011,
24'b110100101011110100101010,
24'b010010001101101100111110,
24'b001011010110001011010110,
24'b000001111101111001011001,
24'b001011010111001011010110,
24'b110010100010111110000001,
24'b001011010110110100101010,
24'b001001101110000010011100,
24'b001011010101001011010110,
24'b110010000011001110001100,
24'b110100101010110100101001,
24'b000000111011110011100000,
24'b001011010110110100101011,
24'b010000011010111111110101,
24'b001011010110001011010110,
24'b111111111010000110000000,
24'b001011010101001011010101,
24'b101111001111010100001110,
24'b110100101010110100101011,
24'b111101110010000100011001,
24'b110100101010110100101010,
24'b000101000111111100001101,
24'b110100101010110100101001,
24'b010100010000101100010110,
24'b001011010110001011010110,
24'b000101011110111010011101,
24'b001011010110001011010111,
24'b111111001110111111111110,
24'b001011010110001011010111,
24'b111000110111000101011010,
24'b001011010110001011010110,
24'b101001101101010011001111,
24'b110100101010110100101010,
24'b110111111111000010011000,
24'b110100101010110100101010,
24'b111101001000110010100101,
24'b001011010101110100101011,
24'b000001000000001001011001,
24'b110100101011110100101010,
24'b000101100010110001010101,
24'b001011010110110100101010,
24'b010001111001111111100000,
24'b001011010111001011010110,
24'b111000110010001101011011,
24'b110100101010110100101010,
24'b001110000000110100000001,
24'b001011010110001011010110,
24'b110101010011000010001011,
24'b001011010101110100101010,
24'b000010101110010001010001,
24'b110100101001110100101010,
24'b001001111000000000100011,
24'b110100101001110100101010,
24'b011001010001101111110100,
24'b001011010110001011010110,
24'b001011001010111110111011,
24'b001011010110001011010111,
24'b000110001111001101000100,
24'b110100101010001011010111,
24'b000010110010110011101000,
24'b001011010110001011010101,
24'b111111100001000001011100,
24'b001011010110001011010101,
24'b111011000111001111010011,
24'b110100101010001011010101,
24'b101110000100110110000101,
24'b001011010110110100101010,
24'b111111111001000100101000,
24'b001011010101110100101001,
24'b010001101111010100100100,
24'b110100101010001011010111,
24'b000100101011000101110110,
24'b110100101011001011010101,
24'b000000010001111110111110,
24'b110100101010001011010110,
24'b111101000000110001101100,
24'b001011010110001011010110,
24'b111001100110001010111010,
24'b110100101010001011010101,
24'b110100110011111100001110,
24'b110100101010001011010110,
24'b100110111100101100001000,
24'b001011010111110100101010,
24'b110111010010111010110010,
24'b001011010110110100101001,
24'b000101111001000001110110,
24'b001011010111001011010101,
24'b101100010110010000001011,
24'b110100101001110100101010,
24'b111000111101111111001101,
24'b110100101010110100101011,
24'b111110100100101110010111,
24'b001011010110110100101010,
24'b001010101000111101010101,
24'b001011010110001011010110,
24'b101111101111001011001101,
24'b110100101010110100101010,
24'b111011010000110001010001,
24'b001011010111110100101010,
24'b111111001100111101110010,
24'b001011010110110100101010,
24'b000010011011000011101001,
24'b001011010110110100101011,
24'b000110100100010000011100,
24'b110100101001110100101011,
24'b010010101110110111100100,
24'b001011010110001011010101,
24'b111001101001001101001010,
24'b110100101010110100101001,
24'b001111001111110101101101,
24'b001011010110001011010110,
24'b110111111100001011101101,
24'b110100101010110100101010,
24'b001110010100110100001111,
24'b001011010110001011010110,
24'b110111101001001001110010,
24'b110100101010110100101010,
24'b001111001000110000110100,
24'b001011010101001011010110,
24'b111111110101111101010100,
24'b001011010110001011010111,
24'b101111100010000010001111,
24'b001011010110110100101011,
24'b111110001110000111011001,
24'b001011010110110100101010,
24'b000101100101010101000010,
24'b110100101010110100101010,
24'b010100100111000011111010,
24'b110100101010001011010110,
24'b000101011011110011010010,
24'b001011010110001011010110,
24'b111101111010000011000011,
24'b001011010110001011010110,
24'b101111000000010011001010,
24'b110100101010110100101010,
24'b111111000001000100000110,
24'b110100101010110100101001,
24'b001101110110111100001111,
24'b110100101010001011010110,
24'b110101001001101100100001,
24'b001011010110110100101011,
24'b000100000001111010100100,
24'b001011010110110100101010,
24'b010100001101111111101001,
24'b001011010101001011010110,
24'b000101101001000011100111,
24'b001011010110001011010110,
24'b111110110011001000011111,
24'b001011010110001011010110,
24'b110001011000010101111110,
24'b110100101001110100101010,
24'b001001110000000100101010,
24'b110100101010001011010101,
24'b110011101101110011100111,
24'b001011010101110100101010,
24'b001010101011000001111101,
24'b001011010110001011010111,
24'b110100000110001001001010,
24'b001011010110110100101010,
24'b001010110001011000000101,
24'b110100101010001011010110,
24'b110011111110001000010111,
24'b110100101010110100101010,
24'b001010010001111010001111,
24'b001011010110001011010110,
24'b110010011010010100010010,
24'b110100101010110100101010,
24'b000001010010001000011011,
24'b110100101011110100101010,
24'b010000110110000100011111,
24'b110100101011001011010110,
24'b000000100001000001100110,
24'b110100101011001011010110,
24'b110000001101111110101111,
24'b110100101010110100101010,
24'b111111110101111010110101,
24'b110100101010110100101010,
24'b001110110001101111000001,
24'b001011010101001011010110,
24'b110111001100001001001001,
24'b110100101010110100101010,
24'b001110011101111011000111,
24'b110100101011001011010111,
24'b111111000111101011100101,
24'b001011010111001011010101,
24'b101110111111111010101010,
24'b001011010110110100101010,
24'b111110011011000001111111,
24'b001011010110110100101010,
24'b001100110000001111111111,
24'b110100101010001011010110,
24'b110011011100111000100011,
24'b001011010110110100101010,
24'b000001010100010000100110,
24'b110100101010110100101010,
24'b001111001001000011010011,
24'b110100101011001011010101,
24'b110101110010111101000101,
24'b110100101010110100101011,
24'b000011110110110000001101,
24'b001011010110110100101010,
24'b010010010110001001101111,
24'b110100101010001011010101,
24'b111010110100111011010111,
24'b110100101010110100101010,
24'b010010100110101011100100,
24'b001011010110001011010110,
24'b000100111000111010100100,
24'b001011010110001011010101,
24'b111101111010000010000110,
24'b001011010110001011010111,
24'b101111001111010001001111,
24'b110100101010110100101010,
24'b111111011000000010001011,
24'b110100101001110100101010,
24'b001110010000111010110101,
24'b110100101010001011010110,
24'b110101100001101100110000,
24'b001011010110110100101010,
24'b000100010000000011111110,
24'b110100101010110100101010,
24'b010011111101101011100000,
24'b001011010110001011010110,
24'b000011111100110111111101,
24'b001011010110001011010111,
24'b110100000111111100010000,
24'b001011010110110100101001,
24'b000100101100111111100000,
24'b001011010101110100101001,
24'b010101101111000011010111,
24'b001011010110001011010111,
24'b000111111111001110101111,
24'b110100101010001011010110,
24'b000010101010110011100110,
24'b001011010110001011010111,
24'b111101010111111111000111,
24'b001011010101001011010110,
24'b101111110001000011011000,
24'b001011010111110100101011,
24'b000001000011000111111001,
24'b001011010110110100101010,
24'b010010000011010100001110,
24'b110100101010001011010101,
24'b000011000101111011001111,
24'b001011010110001011010110,
24'b110100111000010000111010,
24'b110100101001110100101001,
24'b001101100011111001101011,
24'b001011010111001011010110,
24'b111000011100010000001010,
24'b110100101011110100101010,
24'b010001101010111001011101,
24'b001011010111001011010110,
24'b000101001110010000011001,
24'b110100101010001011010101,
24'b111111110101111010011000,
24'b001011010110001011010110,
24'b110011111101010010111010,
24'b110100101011110100101001,
24'b001111000010000101110100,
24'b110100101010001011010111,
24'b000011101000111111101010,
24'b110100101010001011010110,
24'b111111110010110010101101,
24'b001011010110001011010110,
24'b111100100010001011100100,
24'b110100101010001011010111,
24'b111000000101110110010001,
24'b001011010110001011010110,
24'b101010110111001110110110,
24'b110100101010110100101010,
24'b111100001000000000111000,
24'b110100101010110100101010,
24'b001100010001110011000011,
24'b001011010101001011010111,
24'b110101110001001100100000,
24'b110100101010110100101010,
24'b001110011000111110100011,
24'b110100101001001011010110,
24'b000001011011110000001111,
24'b001011010110001011010101,
24'b111011010111001000010000,
24'b110100101010001011010101,
24'b101110011100110001110010,
24'b001011010110110100101010,
24'b000111001010001000000000,
24'b110100101010001011010110,
24'b110001011001101111100010,
24'b001011010110110100101010,
24'b001000100110111100011110,
24'b001011010110001011010111,
24'b110010001100000001101110,
24'b001011010110110100101010,
24'b001000111010000111000100,
24'b001011010110001011010110,
24'b110001100000010100010100,
24'b110100101001110100101010,
24'b000000111010111100100101,
24'b001011010111110100101001,
24'b010001011010010100101111,
24'b110100101010001011010101,
24'b000011000000001000000000,
24'b110100101010001011010110,
24'b111100001000000011011110,
24'b110100101010001011010110,
24'b101101111110000000000011,
24'b110100101010110100101010,
24'b111111001000111100100001,
24'b110100101010110100101010,
24'b010000011001110111100100,
24'b110100101010001011010110,
24'b000010101110101001011101,
24'b001011010110001011010110,
24'b111101010100111000111000,
24'b001011010110001011010110,
24'b110111110101000000000101,
24'b001011010101001011010110,
24'b101001110101001101011111,
24'b110100101001110100101010,
24'b111010011001110100010000,
24'b001011010111110100101010,
24'b001001101111000010110110,
24'b001011010111001011010110,
24'b110010000111010010100111,
24'b110100101001110100101011,
24'b001000011011000010111001,
24'b110100101001001011010111,
24'b110001011000110100010100,
24'b001011010110110100101010,
24'b000111100000001101011000,
24'b110100101010001011011000,
24'b101111010100111111001001,
24'b110100101010110100101001,
24'b111101101001110000100111,
24'b001011010110110100101010,
24'b001011101100001000010000,
24'b110100101011001011010110,
24'b110010100000110000110010,
24'b001011010111110100101010,
24'b000000111000111111100010,
24'b001011010110110100101001,
24'b010000010101001110000000,
24'b110100101010001011010111,
24'b000000001000110101001111,
24'b001011010111001011010101,
24'b110000101110000100010000,
24'b001011010110110100101010,
24'b000111110000010100101111,
24'b110100101010001011010110,
24'b101111101010000110110010,
24'b110100101001110100101010,
24'b111101001010000001100101,
24'b110100101010110100101010,
24'b000100000001111101010110,
24'b110100101010110100101010,
24'b010010100101111000000000,
24'b110100101001001011010110,
24'b000010010100101001100011,
24'b001011010110001011010110,
24'b110011001111111000100101,
24'b001011010110110100101010,
24'b001011001001111110110010,
24'b001011010111001011010110,
24'b110101010011000100110101,
24'b001011010110110100101010,
24'b001101101011010011001111,
24'b110100101010001011010110,
24'b000000001010000011000001,
24'b110100101010001011010110,
24'b111001000110110100000000,
24'b001011010110001011010110,
24'b101010000010001100000001,
24'b110100101010110100101010,
24'b111000111011110110010010,
24'b001011010110110100101010,
24'b111111110100001110101011,
24'b110100101001110100101010,
24'b001101001001000000100111,
24'b110100101010001011010110,
24'b110100100010110010111000,
24'b001011010110110100101010,
24'b001010000010001100101100,
24'b110100101010001011010110,
24'b110001101001111111110111,
24'b110100101010110100101010,
24'b111111111011111001011001,
24'b110100101010110100101010,
24'b001110010101101011001001,
24'b001011010110001011010110,
24'b110110011011111011110101,
24'b001011010110110100101001,
24'b001101011101001100000010,
24'b110100101010001011010111,
24'b111101110101111011110011,
24'b110100101010001011010110,
24'b101101010000101011000111,
24'b001011010110110100101011,
24'b111011100001111001010101,
24'b001011010111110100101010,
24'b000010001000111111110111,
24'b001011010110110100101010,
24'b001111010110001100111000,
24'b110100101011001011010110,
24'b110110110011110011111110,
24'b001011010110110100101010,
24'b001100101001001001000100,
24'b110100101010001011010111,
24'b110101011000101111111110,
24'b001011010110110100101010,
24'b001011100011111100100100,
24'b001011010110001011010110,
24'b110100000000000001111100,
24'b001011010110110100101011,
24'b000110011011001010110010,
24'b000000000001000000000000,
24'b000010001100000100101100,
24'b000000000000000000000000,
24'b000001011100000011001000,
24'b000000000000000000000000,
24'b000001000110000010011000,
24'b000000000000000000000000,
24'b000000111010000001111011,
24'b000000000000000000000000,
24'b000000110001000001100111,
24'b000000000000000000000000,
24'b000000101011000001011000,
24'b000000000000000000000000,
24'b000000100111000001001101,
24'b000000000001000000000000,
24'b000000100011000001000110,
24'b000000000000000000000000,
24'b000000100000000000111111,
24'b000000000000000000000000,
24'b000000011101000000111010,
24'b000000000000000000000000,
24'b000000011011000000110101,
24'b000000000000000000000000,
24'b000000011001000000110001,
24'b000000000000111111111111,
24'b000000011000000000101110,
24'b000000000000000000000000,
24'b000000010111000000101011,
24'b000000000001000000000000,
24'b000000010101000000101001,
24'b000000000000000000000001,
24'b000000010100000000100111,
24'b000000000000000000000001,
24'b000000010010000000100110,
24'b111111111111000000000000,
24'b000000010001000000100011,
24'b000000000000111111111111,
24'b000000010010000000100010,
24'b111111111111000000000000,
24'b000000010000000000100000,
24'b000000000000000000000000,
24'b000000010000000000011111,
24'b000000000000000000000001,
24'b000000001110000000011110,
24'b000000000000000000000000,
24'b000000001110000000011101,
24'b000000000000000000000000,
24'b000000001110000000011100,
24'b000000000000000000000000,
24'b000000001101000000011011,
24'b000000000000000000000000,
24'b000000001100000000011010,
24'b000000000001000000000000,
24'b000000001100000000011010,
24'b000000000000111111111111,
24'b000000001100000000011010,
24'b111111111111000000000000,
24'b000000001100000000011001,
24'b111111111111000000000000,
24'b000000001100000000011000,
24'b000000000000000000000001,
24'b000000001010000000010111,
24'b000000000000111111111111,
24'b000000001011000000010111,
24'b000000000001000000000000,
24'b000000001011000000010111,
24'b111111111111000000000000,
24'b000000001010000000010110,
24'b000000000000000000000000,
24'b000000001011000000010101,
24'b000000000000000000000000,
24'b000000001010000000010101,
24'b000000000000000000000000,
24'b000000001010000000010100,
24'b000000000000000000000000,
24'b000000001001000000010101,
24'b000000000000000000000000,
24'b000000001010000000010100,
24'b000000000000000000000000,
24'b000000001010000000010100,
24'b000000000000000000000001,
24'b000000001001000000010100,
24'b000000000000000000000000,
24'b000000001001000000010011,
24'b000000000000000000000000,
24'b000000001001000000010011,
24'b000000000000000000000000,
24'b000000001001000000010011,
24'b111111111111000000000000,
24'b000000001001000000010010,
24'b000000000000000000000000,
24'b000000001001000000010010,
24'b000000000000000000000000,
24'b000000001000000000010010,
24'b000000000000000000000000,
24'b000000001000000000010001,
24'b000000000000000000000000,
24'b000000001001000000010001,
24'b000000000000000000000001,
24'b000000000111000000010001,
24'b000000000000000000000000,
24'b000000000111000000010001,
24'b000000000000111111111111,
24'b000000001000000000010001,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000001,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000000111000000001111,
24'b000000000000111111111111,
24'b000000000111000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b111111111111000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000000111000000001111,
24'b000000000000000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000001,
24'b000000000111000000001110,
24'b000000000000000000000000,
24'b000000000111000000001110,
24'b000000000000000000000000,
24'b000000000111000000001110,
24'b000000000000000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000000111000000001110,
24'b111111111111000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000000111000000001101,
24'b000000000000000000000000,
24'b000000001000000000001101,
24'b000000000000000000000000,
24'b000000000111000000001101,
24'b111111111111111111111111,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000001000000000001101,
24'b111111111111000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000001000000000001101,
24'b111111111111000000000001,
24'b000000000111000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000001,
24'b000000000111000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000000111000000001100,
24'b000000000001000000000000,
24'b000000001000000000001101,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000000111000000001100,
24'b111111111111000000000000,
24'b000000000111000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b111111111111000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000000111000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000111111111111,
24'b000000001000000000001011,
24'b000000000001000000000001,
24'b000000001000000000001100,
24'b111111111111000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000111111111111,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000111111111111,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000111111111111,
24'b000000001000000000001010,
24'b000000000000111111111111,
24'b000000001001000000001010,
24'b000000000001000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000001000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000001,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000001,
24'b000000001000000000001010,
24'b111111111111000000000000,
24'b000000001001000000001010,
24'b111111111111000000000000,
24'b000000001000000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b111111111111000000000000,
24'b000000001010000000001001,
24'b000000000000000000000001,
24'b000000001000000000001001,
24'b000000000000111111111111,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001010000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000001000000000001,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000111111111111,
24'b000000001001000000001001,
24'b111111111111111111111111,
24'b000000001001000000001001,
24'b111111111111111111111111,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b111111111111000000000001,
24'b000000001001000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000001,
24'b000000001010000000001000,
24'b111111111111000000000000,
24'b000000001010000000000111,
24'b000000000001000000000000,
24'b000000001010000000001000,
24'b111111111111000000000000,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000001,
24'b000000001001000000000111,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b000000000001000000000001,
24'b000000001001000000001000,
24'b111111111111111111111111,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000111111111111,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001011000000001000,
24'b111111111111000000000000,
24'b000000001010000000000110,
24'b000000000001000000000000,
24'b000000001011000000001000,
24'b111111111111000000000001,
24'b000000001010000000000111,
24'b000000000000111111111111,
24'b000000001011000000000111,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b111111111111000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b000000000000111111111111,
24'b000000001011000000000111,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000001000000000000,
24'b000000001011000000000111,
24'b000000000000000000000001,
24'b000000001011000000000111,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b111111111111000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b111111111111111111111111,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000001000000000001,
24'b0_00000001010000000000111,
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b111111111111000000000000, 
24'b000000001010000000000101, 
24'b111111111111000000000001, 
24'b000000001001000000000101, 
24'b000000000000000000000000, 
24'b000000001001000000000101, 
24'b000000000000000000000000, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001010000000000101, 
24'b111111111111000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000111111111111, 
24'b000000001011000000000101, 
24'b000000000000000000000001, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001011000000000101, 
24'b111111111111000000000001, 
24'b000000001001000000000100, 
24'b000000000001000000000000, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001001000000000100, 
24'b000000000000111111111111, 
24'b000000001010000000000100, 
24'b000000000001000000000000, 
24'b000000001011000000000101, 
24'b000000000001000000000001, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001010000000000101, 
24'b000000000000111111111111, 
24'b000000001011000000000101, 
24'b000000000000000000000000, 
24'b000000001010000000000101, 
24'b111111111111000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000001000000000000, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000111111111111, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000101, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000111111111111, 
24'b000000001011000000000011, 
24'b000000000000000000000001, 
24'b000000001010000000000100, 
24'b000000000000111111111111, 
24'b000000001011000000000100, 
24'b000000000001000000000000, 
24'b000000001011000000000101, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000001000000000000, 
24'b000000001010000000000101, 
24'b000000000000111111111111, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000101, 
24'b111111111111000000000000, 
24'b000000001011000000000100, 
24'b111111111111000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000000000000000001, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000001, 
24'b000000001011000000000100, 
24'b111111111111000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000111111111111, 
24'b000000001100000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000111111111111, 
24'b000000001100000000000100, 
24'b111111111111000000000000, 
24'b000000001100000000000011, 
24'b111111111111000000000000, 
24'b000000001011000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b111111111111000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b111111111111000000000000, 
24'b000000001011000000000010, 
24'b000000000000111111111111, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001101000000000010, 
24'b000000000001000000000001, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b111111111111000000000000, 
24'b000000001100000000000001, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000001, 
24'b000000001011000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b111111111111000000000000, 
24'b000000001100000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001100000000000001, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001101000000000010, 
24'b000000000000000000000000, 
24'b000000001100000000000010, 
24'b000000000000000000000000, 
24'b000000001101000000000010, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000010, 
24'b000000000000000000000001, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001100000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000001000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000001, 
24'b000000001100000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000001000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001110000000000010, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b111111111111000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b111111111111000000000000, 
24'b000000001110000000000000, 
24'b000000000000000000000000, 
24'b000000001110000000000000, 
24'b000000000000000000000000, 
24'b000000001110000000000000, 
24'b000000000001000000000000, 
24'b000000001101000000000001, 
24'b000000000000111111111111, 
24'b000000001110000000000001, 
24'b000000000000000000000000, 
24'b000000001101000000000001, 
24'b000000000000000000000000, 
24'b000000001110000000000001, 
24'b111111111111000000000000, 
24'b000000001110000000000000, 
24'b000000000001000000000000, 
24'b000000001110000000000001, 
24'b000000000000000000000000, 
24'b000000001110000000000000, 
24'b000000000000000000000000, 
24'b000000001111000000000000, 
24'b000000000000000000000000, 
24'b000000001111000000000000, 
24'b000000000000000000000001, 
24'b000000001110000000000001, 
24'b111111111111000000000000, 
24'b000000001110000000000000, 
24'b000000000000000000000000, 
24'b000000001111000000000000, 
24'b000000000000000000000000, 
24'b000000001111000000000000, 
24'b000000000000000000000001, 
24'b000000001110111111111111, 
24'b000000000001000000000001, 
24'b000000001110000000000001, 
24'b111111111111000000000000, 
24'b000000001110000000000000, 
24'b000000000000111111111111, 
24'b000000001111000000000000, 
24'b111111111111000000000000, 
24'b000000001111111111111111, 
24'b000000000001000000000000, 
24'b000000001111000000000000, 
24'b000000000000000000000000, 
24'b000000001111000000000000, 
24'b000000000000000000000001, 
24'b000000001111000000000000, 
24'b000000000000000000000000, 
24'b000000001111111111111111, 
24'b000000000000000000000001, 
24'b000000001110111111111111, 
24'b000000000000000000000000, 
24'b000000001111111111111111, 
24'b000000000000000000000000, 
24'b000000001111111111111111, 
24'b000000000000000000000000, 
24'b000000001111111111111111, 
24'b000000000000000000000000, 
24'b000000001111111111111111, 
24'b000000000001000000000000, 
24'b000000010000000000000000, 
24'b000000000000000000000000, 
24'b000000001111111111111111, 
24'b000000000000000000000000, 
24'b000000001111111111111111, 
24'b000000000000111111111111, 
24'b000000010000111111111111, 
24'b000000000000000000000000, 
24'b000000010000111111111111, 
24'b000000000000000000000000, 
24'b000000010000111111111111, 
24'b000000000000000000000000, 
24'b000000010000111111111111, 
24'b111111111111000000000000, 
24'b000000010000111111111110, 
24'b000000000000000000000000, 
24'b000000010000111111111110, 
24'b000000000000000000000000, 
24'b000000010000111111111111, 
24'b000000000000000000000001, 
24'b000000010000111111111111, 
24'b111111111111000000000001, 
24'b000000010000111111111110, 
24'b000000000000000000000000, 
24'b000000010000111111111110, 
24'b000000000000000000000000, 
24'b000000010000111111111110, 
24'b000000000000000000000000, 
24'b000000010000111111111110, 
24'b000000000000000000000000, 
24'b000000010000111111111110, 
24'b000000000000111111111111, 
24'b000000010001111111111110, 
24'b000000000000000000000000, 
24'b000000010001111111111110, 
24'b111111111111000000000000, 
24'b000000010001111111111110, 
24'b111111111111000000000000, 
24'b000000010001111111111101, 
24'b000000000000000000000000, 
24'b000000010001111111111101, 
24'b000000000000000000000000, 
24'b000000010001111111111101, 
24'b000000000001000000000000, 
24'b000000010010111111111110, 
24'b000000000001000000000000, 
24'b000000010010111111111110, 
24'b000000000000000000000000, 
24'b000000010010111111111110, 
24'b000000000000000000000001, 
24'b000000010001111111111101, 
24'b000000000000000000000000, 
24'b000000010010111111111101, 
24'b000000000000000000000000, 
24'b000000010010111111111110, 
24'b000000000000000000000001, 
24'b000000010010111111111101, 
24'b000000000000000000000000, 
24'b000000010011111111111101, 
24'b000000000000000000000000, 
24'b000000010010111111111100, 
24'b000000000001000000000000, 
24'b000000010011111111111101, 
24'b000000000000000000000000, 
24'b000000010011111111111101, 
24'b000000000000000000000000, 
24'b000000010100111111111101, 
24'b000000000000000000000001, 
24'b000000010011111111111101, 
24'b000000000000000000000001, 
24'b000000010010111111111101, 
24'b000000000000000000000000, 
24'b000000010011111111111101, 
24'b000000000000000000000000, 
24'b000000010011111111111101, 
24'b000000000000000000000000, 
24'b000000010011111111111100, 
24'b000000000000000000000000, 
24'b000000010100111111111100, 
24'b000000000000000000000000, 
24'b000000010100111111111101, 
24'b000000000000000000000000, 
24'b000000010100111111111100, 
24'b000000000000000000000000, 
24'b000000010100111111111101, 
24'b000000000000000000000000, 
24'b000000010100111111111100, 
24'b000000000000000000000000, 
24'b000000010101111111111100, 
24'b000000000000000000000001, 
24'b000000010100111111111100, 
24'b000000000000000000000000, 
24'b000000010100111111111011, 
24'b000000000000111111111111, 
24'b000000010110111111111100, 
24'b111111111111000000000000, 
24'b000000010110111111111011, 
24'b000000000000000000000000, 
24'b000000010110111111111011, 
24'b000000000000000000000000, 
24'b000000010110111111111011, 
24'b000000000000000000000000, 
24'b000000010110111111111011, 
24'b000000000000000000000000, 
24'b000000010110111111111011, 
24'b000000000000000000000000, 
24'b000000010111111111111011, 
24'b111111111111000000000000, 
24'b000000010111111111111011, 
24'b000000000000000000000000, 
24'b000000010111111111111011, 
24'b000000000000000000000000, 
24'b000000010111111111111011, 
24'b000000000000000000000000, 
24'b000000010111111111111011, 
24'b000000000000111111111111, 
24'b000000011000111111111010, 
24'b000000000000000000000000, 
24'b000000011000111111111010, 
24'b000000000000000000000000, 
24'b000000011000111111111010, 
24'b000000000000000000000000, 
24'b000000011001111111111010, 
24'b000000000000000000000000, 
24'b000000011001111111111010, 
24'b000000000000000000000000, 
24'b000000011001111111111010, 
24'b000000000000000000000000, 
24'b000000011010111111111010, 
24'b000000000000000000000000, 
24'b000000011001111111111001, 
24'b000000000000000000000000, 
24'b000000011010111111111010, 
24'b000000000000000000000000, 
24'b000000011011111111111001, 
24'b000000000000000000000000, 
24'b000000011011111111111001, 
24'b000000000000000000000000, 
24'b000000011011111111111000, 
24'b000000000001000000000000, 
24'b000000011100111111111001, 
24'b000000000001000000000000, 
24'b000000011100111111111001, 
24'b000000000000000000000001, 
24'b000000011100111111111001, 
24'b000000000000000000000000, 
24'b000000011100111111111001, 
24'b000000000001000000000000, 
24'b000000011101111111111010, 
24'b111111111111000000000000, 
24'b000000011101111111111000, 
24'b000000000000111111111111, 
24'b000000011111111111111000, 
24'b000000000000000000000000, 
24'b000000011111111111111000, 
24'b000000000000000000000000, 
24'b000000011111111111111000, 
24'b000000000000000000000000, 
24'b000000100000111111111000, 
24'b000000000000000000000000, 
24'b000000100000111111111000, 
24'b000000000000000000000000, 
24'b000000100001111111111000, 
24'b000000000000111111111111, 
24'b000000100011111111111000, 
24'b000000000000000000000001, 
24'b000000100010111111110111, 
24'b000000000001000000000001, 
24'b000000100011111111110111, 
24'b000000000001000000000000, 
24'b000000100011111111111000, 
24'b000000000000000000000000, 
24'b000000100100111111110111, 
24'b000000000000000000000000, 
24'b000000100100111111111000, 
24'b111111111111000000000000, 
24'b000000100101111111110111, 
24'b000000000000000000000000, 
24'b000000100111111111110110, 
24'b000000000000000000000001, 
24'b000000100110111111110111, 
24'b111111111111111111111111, 
24'b000000101000111111110101, 
24'b000000000000000000000000, 
24'b000000101001111111110110, 
24'b000000000000111111111111, 
24'b000000101011111111110101, 
24'b000000000000000000000000, 
24'b000000101100111111110101, 
24'b000000000000000000000000, 
24'b000000101101111111110101, 
24'b000000000000000000000001, 
24'b000000101101111111110101, 
24'b000000000000000000000000, 
24'b000000101111111111110101, 
24'b000000000000000000000000, 
24'b000000110001111111110100, 
24'b000000000001000000000000, 
24'b000000110011111111110101, 
24'b000000000000000000000000, 
24'b000000110101111111110011, 
24'b000000000001000000000000, 
24'b000000110110111111110100, 
24'b000000000000000000000001, 
24'b000000110111111111110100, 
24'b000000000000000000000000, 
24'b000000111010111111110011, 
24'b000000000001000000000000, 
24'b000000111101111111110011, 
24'b000000000000000000000001, 
24'b000000111111111111110010, 
24'b000000000000000000000001, 
24'b000001000001111111110010, 
24'b111111111111000000000000, 
24'b000001000101111111110001, 
24'b000000000000000000000001, 
24'b000001000111111111101111, 
24'b000000000000111111111111, 
24'b000001001100111111110000, 
24'b111111111111000000000000, 
24'b000001010000111111101101, 
24'b000000000000111111111111, 
24'b000001010101111111101011, 
24'b000000000000111111111111, 
24'b000001011011111111101010, 
24'b000000000000000000000000, 
24'b000001100000111111100111, 
24'b000000000000111111111111, 
24'b000001101000111111100100, 
24'b000000000000111111111111, 
24'b000001110001111111011111, 
24'b000000000001000000000001, 
24'b000001111001111111011001, 
24'b000000000001000000000000, 
24'b000010000100111111001111, 
24'b000000000000000000000000, 
24'b000010010001111110111101, 
24'b000000000000000000000001, 
24'b000010011011111110011110, 
24'b111111111111000000000000, 
24'b000010011001111101010010, 
24'b000000000000000000000000, 
24'b111111010101110111110111, 
24'b001011010111110100101000, 
24'b010100001101000010010011, 
24'b001011011000001011010111, 
24'b000110111001010000001110, 
24'b110100101000001011011000, 
24'b000001000110110111111111, 
24'b001011010111001011010111, 
24'b110101000010001110010000, 
24'b110100101000110100101001, 
24'b010000000010110111011100, 
24'b001011010111001011010111, 
24'b000100101000001110011001, 
24'b110100101000001011010111, 
24'b000000110111111000010001, 
24'b001011010111001011011000, 
24'b111101110110010000100110, 
24'b110100101001001011011000, 
24'b111010000000000010100011, 
24'b110100101001001011011000, 
24'b101110011001110100111100, 
24'b001011010111110100101000, 
24'b001001000001001111000110, 
24'b110100101000001011011000, 
24'b111011110011000010111000, 
24'b110100101000001011011000, 
24'b101110010000111101111111, 
24'b110100101001110100101001, 
24'b000111101110111000101110, 
24'b110100101001001011010111, 
24'b111001001111101010101011, 
24'b001011010111001011010111, 
24'b101001001101111010100011, 
24'b001011010111110100101000, 
24'b110111101011000010110000, 
24'b001011010111110100101000, 
24'b111101100100010010100110, 
24'b110100101001110100101000, 
24'b000011010111000100011111, 
24'b110100101001110100101000, 
24'b010001011111111111000101, 
24'b110100101001001011010111, 
24'b000000101100111010000000, 
24'b110100101000001011011000, 
24'b110000001111101101011110, 
24'b001011011000110100101000, 
24'b000000000001000111001001, 
24'b110100101001110100101001, 
24'b001111010010111000100110, 
24'b110100101010001011011000, 
24'b111000001100101000011110, 
24'b001011010110110100101000, 
24'b010000100001110110101101, 
24'b001011011000001011010111, 
24'b000011100001111100010101, 
24'b001011011000001011010111, 
24'b111110001100000001100111, 
24'b001011010111001011010111, 
24'b111000100100001110011100, 
24'b110100101001001011010111, 
24'b101010001101110101101111, 
24'b001011010111110100101000, 
24'b111001110000001011101000, 
24'b110100101001110100101000, 
24'b000001100000110100011110, 
24'b001011011000110100101001, 
24'b010000100010001010111110, 
24'b110100101001001011011000, 
24'b000000100000110100001001, 
24'b001011010111001011011000, 
24'b110001011111001010111001, 
24'b110100101001110100101000, 
24'b001001011011110100011110, 
24'b001011010111001011011000, 
24'b110011001101001100010100, 
24'b110100101000110100101001, 
24'b001010011001111101100000, 
24'b110100101000001011010111, 
24'b110100010101101110100100, 
24'b001011010111110100101001, 
24'b001100101011000101111011, 
24'b110100101001001011011000, 
24'b111111000011101110000110, 
24'b001011010111001011010111, 
24'b110111111000111100011101, 
24'b001011011000001011010111, 
24'b101000100111001010011101, 
24'b110100101000110100101000, 
24'b110111001001110000111010, 
24'b001011011000110100101001, 
24'b111100110111111110110010, 
24'b001011010111110100101001, 
24'b000010011001001100110011, 
24'b110100101001110100101001, 
24'b010000001010110100010000, 
24'b001011011000001011011000, 
24'b111110110011001001110101, 
24'b110100101000001011011000, 
24'b101101011111110001011100, 
24'b001011011000110100101000, 
24'b111011011010111111111111, 
24'b001011011000110100101000, 
24'b000001101100001111011000, 
24'b110100101000110100101001, 
24'b001110011101111110111101, 
24'b110100101001001011010111, 
24'b110100101101101111001100, 
24'b001011010111110100101001, 
24'b000010110101000101110110, 
24'b110100101000110100101000, 
24'b010010001011101101000100, 
24'b001011010111001011011000, 
24'b000001111000111001100010, 
24'b001011011000001011011000, 
24'b110010011010111110001010, 
24'b001011010111110100101001, 
24'b001001101001000010100101, 
24'b001011010111001011010111, 
24'b110001111011001110011000, 
24'b110100101000110100101001, 
24'b000000110011110011101001, 
24'b001011010111110100101000, 
24'b010000010111111111111110, 
24'b001011011000001011011000, 
24'b111111110101000110001011, 
24'b001011010111001011011000, 
24'b101111000110010100011011, 
24'b110100101001110100101000, 
24'b111101101101000100100101, 
24'b110100101000110100101000, 
24'b000101000011111100010111, 
24'b110100101000110100101001, 
24'b010100001100101100011111, 
24'b001011010111001011010111, 
24'b000101011001111010101000, 
24'b001011010111001011011000, 
24'b111111001001000000001000, 
24'b001011011000001011011000, 
24'b111000110001000101100110, 
24'b001011011000001011010111, 
24'b101001100101010011011100, 
24'b110100101001110100101001, 
24'b110111110111000010100100, 
24'b110100101000110100101000, 
24'b111101000010110010101110, 
24'b001011011000110100101000, 
24'b000000111100001001100111, 
24'b110100101000110100101001, 
24'b000101011111110001011101, 
24'b001011011000110100101001, 
24'b010001110111111111101011, 
24'b001011011000001011011000, 
24'b111000101100001101101000, 
24'b110100101000110100101000, 
24'b001101111101110100001010, 
24'b001011011000001011011000, 
24'b110101001110000010010101, 
24'b001011011000110100101001, 
24'b000010101010010001011111, 
24'b110100101001110100101001, 
24'b001001110100000000101111, 
24'b110100101001110100101000, 
24'b011001001111101111111111, 
24'b001011011000001011010111, 
24'b001011000110111111001000, 
24'b001011010111001011011000, 
24'b000110001010001101010010, 
24'b110100101000001011010111, 
24'b000010101111110011110011, 
24'b001011010111001011010111, 
24'b111111011100000001101000, 
24'b001011011000001011010111, 
24'b111011000001001111100001, 
24'b110100101001001011010111, 
24'b101101111101110110010000, 
24'b001011010111110100101000, 
24'b111111110100000100110101, 
24'b001011010111110100101001, 
24'b010001101011010100110011, 
24'b110100101001001011010110, 
24'b000100100111000110000100, 
24'b110100101001001011010111, 
24'b000000001101111111001011, 
24'b110100101000001011010110, 
24'b111100111100110001110111, 
24'b001011010111001011011000, 
24'b111001100010001011001000, 
24'b110100101000001011011000, 
24'b110100101101111100011010, 
24'b110100101000001011011000, 
24'b100110110100101100010010, 
24'b001011011000110100101001, 
24'b110111001100111010111110, 
24'b001011011000110100101001, 
24'b000101110101000010000011, 
24'b001011010111001011010111, 
24'b101100001110010000011000, 
24'b110100101001110100101001, 
24'b111000110101111111011010, 
24'b110100101001110100101001, 
24'b111110011111101110100001, 
24'b001011011000110100101000, 
24'b001010100100111101100001, 
24'b001011010111001011011000, 
24'b101111101000001011011010, 
24'b110100101010110100101001, 
24'b111011001011110001011101, 
24'b001011011000110100101000, 
24'b111111000110111101111111, 
24'b001011010111110100101000, 
24'b000010010110000011110110, 
24'b001011011000110100101001, 
24'b000110100000010000101011, 
24'b110100101001110100101001, 
24'b010010101100110111110001, 
24'b001011010111001011010111, 
24'b111001100011001101011001, 
24'b110100101001110100101000, 
24'b001111001101110101111010, 
24'b001011010111001011011001, 
24'b110111110101001011111011, 
24'b110100101001110100101000, 
24'b001110010001110100011011, 
24'b001011010111001011011000, 
24'b110111100010001010000001, 
24'b110100101000110100101000, 
24'b001111000101110000111111, 
24'b001011011000001011011000, 
24'b111111101111111101100010, 
24'b001011010111001011010111, 
24'b101111011011000010011101, 
24'b001011011000110100101001, 
24'b111110001010000111101000, 
24'b001011011000110100101001, 
24'b000101100000010101010011, 
24'b110100101000110100100111, 
24'b010100100101000100001000, 
24'b110100101001001011010111, 
24'b000101011000110011011111, 
24'b001011011000001011011000, 
24'b111101110101000011010010, 
24'b001011010111001011010111, 
24'b101110111010010011011010, 
24'b110100101001110100101001, 
24'b111110111100000100010101, 
24'b110100101000110100101001, 
24'b001101110010111100011101, 
24'b110100101001001011011000, 
24'b110101000010101100101110, 
24'b001011010111110100101001, 
24'b000011111100111010110010, 
24'b001011010111110100101000, 
24'b010100001011111111110111, 
24'b001011010111001011011000, 
24'b000101100100000011110110, 
24'b001011010111001011010111, 
24'b111110101110001000101110, 
24'b001011010111001011011000, 
24'b110001010001010110010000, 
24'b110100100111110100101000, 
24'b001001101100000100111001, 
24'b110100101001001011010111, 
24'b110011100101110011110100, 
24'b001011010111110100101000, 
24'b001010100111000010001101, 
24'b001011010111001011010111, 
24'b110100000000001001011011, 
24'b001011011000110100101001, 
24'b001010101110011000011000, 
24'b110100101000001011010111, 
24'b110011110111001000101000, 
24'b110100101000110100101000, 
24'b001010001110111010011110, 
24'b001011010111001011011000, 
24'b110010010011010100100100, 
24'b110100101001110100101000, 
24'b000001001101001000101100, 
24'b110100101001110100101001, 
24'b010000110100000100101111, 
24'b110100101001001011011000, 
24'b000000011100000001110111, 
24'b110100101001001011011000, 
24'b110000000101111110111111, 
24'b110100101000110100101000, 
24'b111111110000111011000011, 
24'b110100101000110100101000, 
24'b001110101110101111001110, 
24'b001011010111001011010111, 
24'b110111000110001001011010, 
24'b110100101001110100101001, 
24'b001110011010111011011000, 
24'b110100101001001011011000, 
24'b111111000010101011110010, 
24'b001011010111001011010111, 
24'b101110110111111010111001, 
24'b001011011000110100101000, 
24'b111110010101000010010000, 
24'b001011010111110100101000, 
24'b001100101101010000010011, 
24'b110100101000001011010111, 
24'b110011010110111000110011, 
24'b001011011000110100101001, 
24'b000001001111010000111011, 
24'b110100100111110100101001, 
24'b001111000110000011100101, 
24'b110100101000001011011000, 
24'b110101101010111101010101, 
24'b110100101000110100101000, 
24'b000011110010110000011011, 
24'b001011011000110100101001, 
24'b010010010100001010000010, 
24'b110100101000001011010111, 
24'b111010101110111011100110, 
24'b110100101001110100101000, 
24'b010010100011101011110010, 
24'b001011010111001011010111, 
24'b000100110011111010110100, 
24'b001011011000001011010111, 
24'b111101110011000010011000, 
24'b001011011000001011010111, 
24'b101111000111010001100011, 
24'b110100101001110100101000, 
24'b111111010010000010011111, 
24'b110100100111110100101000, 
24'b001110001011111011000111, 
24'b110100101000001011010111, 
24'b110101011010101101000000, 
24'b001011010111110100101000, 
24'b000100001011000100010001, 
24'b110100101001110100101000, 
24'b010011111010101011110000, 
24'b001011010111001011010111, 
24'b000011110110111000001111, 
24'b001011010111001011010111, 
24'b110100000010111100100010, 
24'b001011010111110100101000, 
24'b000100100111111111110011, 
24'b001011011000110100101000, 
24'b010101101100000011101100, 
24'b001011011000001011010111, 
24'b000111111011001111000101, 
24'b110100101000001011011000, 
24'b000010100100110011111000, 
24'b001011010111001011010111, 
24'b111101010010111111011011, 
24'b001011010111001011010111, 
24'b101111101010000011101101, 
24'b001011011000110100101000, 
24'b000000111110001000001111, 
24'b001011010111110100101000, 
24'b010010000010010100100110, 
24'b110100101000001011011000, 
24'b000011000000111011100010, 
24'b001011011000001011011000, 
24'b110100110000010001010010, 
24'b110100101001110100101001, 
24'b001101011110111010000001, 
24'b001011011000001011011000, 
24'b111000010101010000100010, 
24'b110100101001110100101001, 
24'b010001100101111001110011, 
24'b001011010110001011010111, 
24'b000101001001010000110000, 
24'b110100101000001011010111, 
24'b111111101110111010101101, 
24'b001011010111001011011001, 
24'b110011110101010011010010, 
24'b110100101001110100101000, 
24'b001110111100000110001100, 
24'b110100101000001011011000, 
24'b000011100010111111111111, 
24'b110100101001001011011000, 
24'b111111101010110011000010, 
24'b001011011000001011010111, 
24'b111100011010001011111110, 
24'b110100101000001011011000, 
24'b110111111110110110100110, 
24'b001011010111001011010111, 
24'b101010101110001111010000, 
24'b110100101001110100101000, 
24'b111100000001000001010000, 
24'b110100101000110100101000, 
24'b001100001100110011011001, 
24'b001011010111001011010111, 
24'b110101101010001100111011, 
24'b110100101000110100101001, 
24'b001110010011111110111100, 
24'b110100101000001011011000, 
24'b000001010100110000100111, 
24'b001011011000001011011000, 
24'b111011001111001000101011, 
24'b110100101000001011010111, 
24'b101110010010110010001010, 
24'b001011011000110100101001, 
24'b000111000011001000011100, 
24'b110100101000001011011000, 
24'b110001001111101111111011, 
24'b001011010111110100101000, 
24'b001000100000111100111000, 
24'b001011010111001011011000, 
24'b110010000011000010001001, 
24'b001011010111110100101010, 
24'b001000110010000111100000, 
24'b001011011000001011010111, 
24'b110001010101010100110100, 
24'b110100101000110100101000, 
24'b000000110011111101000010, 
24'b001011010111110100101000, 
24'b010001010100010101001101, 
24'b110100101001001011010111, 
24'b000010111000001000011110, 
24'b110100101001001011010111, 
24'b111011111111000011111100, 
24'b110100101000001011011000, 
24'b101101110011000000100001, 
24'b110100101000110100101000, 
24'b111110111111111101000000, 
24'b110100101000110100101001, 
24'b010000010010111000000010, 
24'b110100101001001011011000, 
24'b000010100101101001111010, 
24'b001011011000001011011000, 
24'b111101001010111001010111, 
24'b001011010111001011010111, 
24'b110111101001000000100101, 
24'b001011011000001011011000, 
24'b101001100111001110000011, 
24'b110100101000110100101000, 
24'b111010001110110100110010, 
24'b001011010111110100101000, 
24'b001001100110000011011000, 
24'b001011011000001011011000, 
24'b110001111010010011001100, 
24'b110100101000110100101001, 
24'b001000010001000011011110, 
24'b110100101000001011011000, 
24'b110001001011110100111000, 
24'b001011010111110100101000, 
24'b000111010110001101111111, 
24'b110100101000001011010111, 
24'b101111001001111111101101, 
24'b110100101001110100101001, 
24'b111101011101110001001011, 
24'b001011010111110100101001, 
24'b001011100010001000110111, 
24'b110100101001001011011000, 
24'b110010010010110001011000, 
24'b001011011000110100101000, 
24'b000000101100000000001010, 
24'b001011011000110100101001, 
24'b010000001010001110101011, 
24'b110100101000001011011000, 
24'b111111111011110101111000, 
24'b001011011000001011010111, 
24'b110000011110000100111101, 
24'b001011010111110100101000, 
24'b000111100011010101011101, 
24'b110100101001001011010111, 
24'b101111011010000111011111, 
24'b110100101010110100101000, 
24'b111100111100000010010101, 
24'b110100101001110100101000, 
24'b000011110011111110000110, 
24'b110100101001110100101000, 
24'b010010011001111000110000, 
24'b110100101000001011011000, 
24'b000010000101101010010011, 
24'b001011010111001011010111, 
24'b110010111101111001011000, 
24'b001011010111110100101001, 
24'b001010111010111111100111, 
24'b001011011000001011011000, 
24'b110101000001000101101101, 
24'b001011010111110100101000, 
24'b001101011100010100001010, 
24'b110100101000001011010111, 
24'b111111111000000011111011, 
24'b110100101000001011010111, 
24'b111000110010110100111011, 
24'b001011010111001011011000, 
24'b101001101010001101000001, 
24'b110100101000110100101000, 
24'b111000100101110111010010, 
24'b001011011000110100101001, 
24'b111111011101001111110001, 
24'b110100101001110100101000, 
24'b001100110010000001110010, 
24'b110100101000001011010111, 
24'b110100000101110100000110, 
24'b001011010111110100101001, 
24'b001001100011001110000110, 
24'b110100101001001011010111, 
24'b110000111110000001100001, 
24'b110100101000110100101010, 
24'b111110110011111011101110, 
24'b110100101001110100101010, 
24'b001001101100110001101111, 
24'b000000000001111111111111, 
24'b001000010011110010011111, 
24'b001011010111001011010111, 
24'b110100100111111110101010, 
24'b001011010111110100101000, 
24'b001100010101001110000111, 
24'b110100101000001011010111, 
24'b111100111010111101100101, 
24'b110100101001001011011000, 
24'b101100010110101100110001, 
24'b001011011000110100101001, 
24'b111010101010111011000000, 
24'b001011011000110100101000, 
24'b000001010000000001100010, 
24'b001011010111110100101000, 
24'b001110011101001110101000, 
24'b110100101000001011011000, 
24'b110101101111110101101100, 
24'b001011011000110100101000, 
24'b001011011111001010111000, 
24'b110100101000001011011000, 
24'b110011111011110001101111, 
24'b001011010111110100101000, 
24'b001001101011111110010010, 
24'b001011010111001011011000, 
24'b110000111110000011001111, 
24'b001011010111110100101001, 
24'b111110001101001000010101, 
24'b001011011000110100101001, 
24'b000100111010010101010101, 
24'b110100101001110100101001, 
24'b010011011111111101001101, 
24'b001011010111001011010111, 
24'b000011111001010100101101, 
24'b110100101001001011011000, 
24'b111011110110000110010001, 
24'b110100101001001011011000, 
24'b101100001100111000011111, 
24'b001011011000110100101001, 
24'b111010101001010010101001, 
24'b110100101000110100101000, 
24'b000001000110000110100110, 
24'b110100101001110100101001, 
24'b001101110001000010010000, 
24'b110100101001001011011000, 
24'b110011100000111110100010, 
24'b110100101001110100101001, 
24'b000000001010111001100100, 
24'b110100101001110100101001, 
24'b000110100011101011100010, 
24'b001011011000110100101001, 
24'b010100110101111011001100, 
24'b001011010111001011010111, 
24'b000100011001000010101111, 
24'b001011010111001011010111, 
24'b110101010010010000110000, 
24'b110100101000110100101001, 
24'b001101111000111000111001, 
24'b001011011000001011011000, 
24'b111110111100001111101010, 
24'b110100101000001011010111, 
24'b101110111100111001100011, 
24'b001011010111110100101000, 
24'b111110100001010001111111, 
24'b110100101000110100101001, 
24'b001100111101000100000010, 
24'b110100101001001011010111, 
24'b110011101100110110011111, 
24'b001011010111110100101000, 
24'b000001101110010000100010, 
24'b110100101001110100101001, 
24'b001111110001000011011010, 
24'b110100101001001011010111, 
24'b110110101011110110100011, 
24'b001011010111110100101000, 
24'b000101011110010001011111, 
24'b110100101001110100101001, 
24'b010101101101000110010011, 
24'b110100101000001011010111, 
24'b000111011100000010111111, 
24'b110100101000001011011000, 
24'b000001101011000000110101, 
24'b110100101000001011010111, 
24'b111100000010111111000001, 
24'b110100101001001011011000, 
24'b101110000010111101010001, 
24'b110100101001110100101000, 
24'b111110111110111011010111, 
24'b110100101001110100101000, 
24'b001111100011111000111100, 
24'b110100101001001011011000, 
24'b111111111001110101001010, 
24'b110100101001001011011000, 
24'b110000110010101001000001, 
24'b001011011000110100101001, 
24'b001000000100000001111000, 
24'b110100101001001011011000, 
24'b110000000000101011000001, 
24'b001011010111110100101000, 
24'b111101100000111010001011, 
24'b001011011000110100101000, 
24'b000100000101001001000001, 
24'b110100101001110100101000, 
24'b010001100011110000111100, 
24'b001011010111001011011000, 
24'b111001010101000110101101, 
24'b110100101001110100101000, 
24'b001111111011101110001001, 
24'b001011011000001011011000, 
24'b111001110100111011011111, 
24'b001011011000110100101001, 
24'b010010101000000010001001, 
24'b001011011000001011011000, 
24'b000110001001010000011010, 
24'b110100101001001011011000, 
24'b000001101101111111100011, 
24'b110100101000001011011000, 
24'b111110010100101110111010, 
24'b001011010111001011011000, 
24'b111010101110111110010101, 
24'b001011010111001011010111, 
24'b110101101000001101000010, 
24'b110100101001001011010111, 
24'b100111010000110100111000, 
24'b001011011001110100101010, 
24'b110110001101001010110010, 
24'b110100101001110100101000, 
24'b111100001110110010101100, 
24'b001011010111110100101001, 
24'b000001111000000001011111, 
24'b001011010111110100101000, 
24'b001111101101010001000101, 
24'b110100101001001011010111, 
24'b111110010110000000110011, 
24'b110100101001001011010111, 
24'b101100111110110000100100, 
24'b001011010111110100101000, 
24'b111010101101000000011001, 
24'b001011011000110100101001, 
24'b000000101011001111101011, 
24'b110100101000110100101010, 
24'b001100110111111000011111, 
24'b001011011000001011011000, 
24'b110010000001010000101001, 
24'b110100101000110100101001, 
24'b111101101000000011001011, 
24'b110100101000110100101000, 
24'b000001100110111100011110, 
24'b110100101001110100101000, 
24'b000100110001101110001111, 
24'b001011010111110100101000, 
24'b001000010000111111000111, 
24'b001011010111110100101001, 
24'b001101010111001111110001, 
24'b110100101001110100101000, 
24'b011011111100000000010101, 
24'b110100101001001011010111, 
24'b001101010111110001100000, 
24'b001011010111001011011000, 
24'b001000001100001001010010, 
24'b110100101000001011011000, 
24'b000100101010110010000110, 
24'b001011011000001011010111, 
24'b000001011010000001101000, 
24'b001011010111001011011000, 
24'b111101010001010001111101, 
24'b110100101000001011011000, 
24'b110001001110000010101101, 
24'b110100101001110100101001, 
24'b001010110001110100101101, 
24'b001011010111001011010111, 
24'b110110000011001110101011, 
24'b110100101001110100101001, 
24'b001111100011000010011000, 
24'b110100101001001011010111, 
24'b000011011000111101011011, 
24'b110100101000001011011000, 
24'b111110110101111000000101, 
24'b110100101001001011010111, 
24'b111010010111101001111110, 
24'b001011010111001011011000, 
24'b101110010111111001110000, 
24'b001011011000110100100111, 
24'b001000110101000001110111, 
24'b001011010111001011011000, 
24'b111100000010010001100011, 
24'b110100101000001011010111, 
24'b110101001100000011001011, 
24'b110100101000001011011000, 
24'b100101111100111101010101, 
24'b110100101000110100101001, 
24'b110100001001110111011101, 
24'b110100101001110100101001, 
24'b111001000011101001000010, 
24'b001011010111110100101001, 
24'b111100010111111001000011, 
24'b001011010111110100100111, 
24'b111111011010000111011011, 
24'b110100101001110100101000, 
24'b000011001101101101100011, 
24'b001011011000110100101000, 
24'b001110101000111001101100, 
24'b001011011000001011011000, 
24'b110011011110111101111101, 
24'b001011011000110100101000, 
24'b111111000111000001010010, 
24'b001011010111110100101000, 
24'b000011100000000100110010, 
24'b001011011000110100101000, 
24'b001000001100001001110101, 
24'b001011011000110100101001, 
24'b010100110100011000000101, 
24'b110100101000001011010111, 
24'b111100010011001000110010, 
24'b110100101000110100101000, 
24'b010011010111000001101110, 
24'b110100101001001011010111, 
24'b000100010010110100011011, 
24'b001011011000001011010111, 
24'b110101011100001101010101, 
24'b110100101000110100101000, 
24'b001101010101111000010000, 
24'b001011010111001011011000, 
24'b110110111101010001101010, 
24'b110100101001110100101000, 
24'b001101101110000101101001, 
24'b110100101000001011010111, 
24'b110110010101000001100111, 
24'b110100101001110100101001, 
24'b000101111110111110101000, 
24'b110100101001110100101001, 
24'b010110111010111011100100, 
24'b110100101001001011010111, 
24'b001001011001110111001010, 
24'b110100101001001011010111, 
24'b000100110001101001111011, 
24'b001011011000001011011000, 
24'b000001011110111011011001, 
24'b001011010111001011010111, 
24'b111110001111001100010011, 
24'b110100101000001011011000, 
24'b111001101111111100110110, 
24'b110100101001001011011000, 
24'b101100011110101101010110, 
24'b001011011000110100101001, 
24'b111101111101111110000101, 
24'b001011010111110100101001, 
24'b001111000010001111000111, 
24'b110100101001001011011000, 
24'b111111111111000001001101, 
24'b110100101001001011010111, 
24'b110001110010111011100011, 
24'b110100101001110100101000, 
24'b001011000001110101101110, 
24'b110100101001001011011000, 
24'b111100100101100111001001, 
24'b001011010111001011010111, 
24'b101101000100110110011001, 
24'b001011010111110100101001, 
24'b111101001001111101101011, 
24'b001011010111110100101000, 
24'b001100011000001100000011, 
24'b110100101010001011011000, 
24'b110100110110111010111010, 
24'b110100101000110100101001, 
24'b001100001000101001011101, 
24'b001011011000001011011000, 
24'b111100100011110110110101, 
24'b001011010111001011010111, 
24'b101011110100111011011111, 
24'b001011011000110100101001, 
24'b111001100101111111001011, 
24'b001011010111110100101000, 
24'b111110100110000011101110, 
24'b001011011000110100101000, 
24'b000010100011010000110111, 
24'b110100101001110100101001, 
24'b000111010010111111000001, 
24'b110100101001110100101000, 
24'b010100000001101101001010, 
24'b001011010111001011010111, 
24'b111011011101111010010000, 
24'b001011011000110100101000, 
24'b010001110100111110110010, 
24'b001011010111001011011000, 
24'b111011100011000010010011, 
24'b001011010111110100101001, 
24'b010100001011000110101010, 
24'b001011010111001011010111, 
24'b000111010010010011000000, 
24'b110100101000001011011000, 
24'b000001100100111010000001, 
24'b001011011000001011011000, 
24'b110101011110001111110101, 
24'b110100101001110100101001, 
24'b010000011101111000101110, 
24'b001011010111001011010111, 
24'b000101000001001111011011, 
24'b110100101000001011011000, 
24'b000001001101111001001000, 
24'b001011011000001011011000, 
24'b111110001011010001010101, 
24'b110100101001001011011001, 
24'b111010010010000011001100, 
24'b110100101001001011011000, 
24'b101110101010110101011111, 
24'b001011010111110100101000, 
24'b001001010000001111100100, 
24'b110100101000001011010111, 
24'b111100000001000011010001, 
24'b110100101000001011011000, 
24'b101110011101111110010110, 
24'b110100101001110100101001, 
24'b000111111011111001000010, 
24'b110100101000001011011000, 
24'b111001011001101010111011, 
24'b001011010111001011010111, 
24'b101001011000111010110001, 
24'b001011011000110100101001, 
24'b110111110100000010111101, 
24'b001011010111110100101001, 
24'b111101101100010010110010, 
24'b110100101000110100101000, 
24'b000011100000000100101000, 
24'b110100101000110100101001, 
24'b010001100110111111001100, 
24'b110100101000001011011000, 
24'b000000110010111010000110, 
24'b110100101000001011011000, 
24'b110000010101101101100011, 
24'b001011011000110100101000, 
24'b000000000110000111001101, 
24'b110100101001110100101000, 
24'b001111011000111000101010, 
24'b110100101001001011011000, 
24'b111000010001101000100000, 
24'b001011010111110100101001, 
24'b010000100101110110110000, 
24'b001011011000001011010111, 
24'b000011100101111100010111, 
24'b001011010111001011011000, 
24'b111110001110000001100111, 
24'b001011011000001011010111, 
24'b111000101000001110011110, 
24'b110100101001001011011000, 
24'b101010010000110101101111, 
24'b001011010111110100101001, 
24'b111001110011001011100111, 
24'b110100101001110100101000, 
24'b000001100010110100011101, 
24'b001011011001110100101000, 
24'b010000100101001010111101, 
24'b110100101001001011011000, 
24'b000000100011110100000111, 
24'b001011010111001011011001, 
24'b110001100001001010111000, 
24'b110100101001110100101000, 
24'b001001011101110100011100, 
24'b001011010111001011011000, 
24'b110011001110001100010010, 
24'b110100101000110100101000, 
24'b001010011010111101011110, 
24'b110100101000001011010111, 
24'b110100010110101110100010, 
24'b001011010111110100101000, 
24'b001100101100000101111001, 
24'b110100101000001011010111, 
24'b111111000110101110000010, 
24'b001011011000001011010111, 
24'b110111111010111100011010, 
24'b001011010111001011011000, 
24'b101000101000001010011010, 
24'b110100101000110100100111, 
24'b110111001010110000110111, 
24'b001011010110110100101001, 
24'b111100111001111110101101, 
24'b001011011000110100101001, 
24'b000010011010001100110000, 
24'b110100101000110100101001, 
24'b010000001010110100001100, 
24'b001011011000001011011000, 
24'b111110110100001001110001, 
24'b110100101000001011011000, 
24'b101101100000110001011000, 
24'b001011011000110100101001, 
24'b111011011010111111111100, 
24'b001011010111110100101001, 
24'b000001101011001111010100, 
24'b110100101000110100101000, 
24'b001110011101111110111001, 
24'b110100101000001011010111, 
24'b110100101101101111001000, 
24'b001011010110110100101001, 
24'b000010110101000101110001, 
24'b110100101001110100101000, 
24'b010010001010101101000000, 
24'b001011011000001011011000, 
24'b000001111000111001011111, 
24'b001011011000001011011000, 
24'b110010011010111110000111, 
24'b001011011000110100101001, 
24'b001001101001000010100010, 
24'b001011010111001011011000, 
24'b110001111011001110010101, 
24'b110100101001110100101000, 
24'b000000110101110011100110, 
24'b001011010111110100101000, 
24'b010000010111111111111011, 
24'b001011011000001011011000, 
24'b111111110100000110001001, 
24'b001011010111001011011000, 
24'b101111000111010100011001, 
24'b110100101000110100101000, 
24'b111101101100000100100010, 
24'b110100101001110100101000, 
24'b000101000011111100010101, 
24'b110100101000110100101000, 
24'b010100001101101100011100, 
24'b001011010111001011011000, 
24'b000101011000111010100101, 
24'b001011011000001011010111, 
24'b111111001000000000001000, 
24'b001011010111001011010111, 
24'b111000110010000101100101, 
24'b001011010111001011010111, 
24'b101001100110010011011011, 
24'b110100101001110100101000, 
24'b110111111001000010100100, 
24'b110100100111110100101000, 
24'b111101000010110010101101, 
24'b001011010111110100101000, 
24'b000000111100001001100111, 
24'b110100101000110100101000, 
24'b000101100000110001011110, 
24'b001011011000110100101001, 
24'b010001111000111111101100, 
24'b001011011000001011010111, 
24'b111000101110001101101000, 
24'b110100101001110100101001, 
24'b001101111111110100001101, 
24'b001011010111001011010111, 
24'b110101001111000010011000, 
24'b001011010111110100101001, 
24'b000010101100010001100001, 
24'b110100101001110100101000, 
24'b001001110111000000110010, 
24'b110100101000110100101000, 
24'b011001010011110000000001, 
24'b001011011000001011011000, 
24'b001011001010111111001011, 
24'b001011011000001011011000, 
24'b000110001111001101010111, 
24'b110100101001001011011000, 
24'b000010110011110011111001, 
24'b001011010111001011011000, 
24'b111111100001000001101111, 
24'b001011011000001011010111, 
24'b111011000111001111101001, 
24'b110100101001001011011000, 
24'b101110000010110110011000, 
24'b001011011000110100101000, 
24'b111111111011000100111111, 
24'b001011010111110100101001, 
24'b010001110100010100111111, 
24'b110100101000001011011000, 
24'b000100110000000110010000, 
24'b110100101000001011011000, 
24'b000000010111111111011000, 
24'b110100101000001011011000, 
24'b111101000110110010000110, 
24'b001011010111001011010111, 
24'b111001101110001011011001, 
24'b110100101000001011011000, 
24'b110100111100111100101101, 
24'b110100101000001011011000, 
24'b100111000101101100100111, 
24'b001011011000110100101001, 
24'b110111100000111011010111, 
24'b001011010111110100101000, 
24'b000110001110000010011101, 
24'b001011011000001011010111, 
24'b101100101011010000111001, 
24'b110100101000110100101001, 
24'b111001011001111111111110, 
24'b110100101001110100101001, 
24'b111111001011101111001101, 
24'b001011010111110100101000, 
24'b001011011110111110010011, 
24'b001011011000001011011000, 
24'b110000110101001100011011, 
24'b110100101001110100101001, 
24'b111100111010110010110001, 
24'b001011011000110100101001, 
24'b000010000100000000000100, 
24'b001011011000110100101001, 
24'b001010110010001010001011, 
24'b000000000000111111111111, 
24'b000100100111000100011111, 
24'b000000000000000000000000, 
24'b000011000000000011001001, 
24'b000000000000000000000000, 
24'b000010001110000010011111, 
24'b000000000000000000000000, 
24'b000001101111000010000111, 
24'b000000000000000000000000, 
24'b000001011011000001110111, 
24'b000000000000000000000000, 
24'b000001001100000001101011, 
24'b000000000000000000000000, 
24'b000001000010000001100001, 
24'b000000000000000000000000, 
24'b000000111001000001011001, 
24'b000000000000000000000000, 
24'b000000110011000001010100, 
24'b000000000000000000000000, 
24'b000000101101000001001111, 
24'b000000000000111111111111, 
24'b000000101001000001001010, 
24'b000000000000111111111111, 
24'b000000100110000001000110, 
24'b000000000000000000000000, 
24'b000000100011000001000011, 
24'b000000000000000000000001, 
24'b000000011111000001000001, 
24'b111111111111000000000000, 
24'b000000011101000000111101, 
24'b000000000001000000000000, 
24'b000000011011000000111100, 
24'b000000000000000000000000, 
24'b000000011001000000111001, 
24'b000000000001000000000000, 
24'b000000011000000000110111, 
24'b000000000001111111111111, 
24'b000000010111000000110110, 
24'b000000000000111111111111, 
24'b000000010110000000110100, 
24'b000000000000000000000000, 
24'b000000010100000000110010, 
24'b000000000000000000000000, 
24'b000000010100000000110001, 
24'b000000000000000000000000, 
24'b000000010011000000101111, 
24'b000000000000000000000001, 
24'b000000010010000000101111, 
24'b111111111111000000000000, 
24'b000000010001000000101011, 
24'b000000000001000000000000, 
24'b000000010001000000101100, 
24'b000000000000000000000000, 
24'b000000010000000000101010, 
24'b000000000000000000000001, 
24'b000000001111000000101010, 
24'b000000000000000000000000, 
24'b000000001110000000101001, 
24'b000000000000111111111111, 
24'b000000001111000000101000, 
24'b000000000000000000000000, 
24'b000000001110000000101000, 
24'b111111111111111111111111, 
24'b000000001111000000100110, 
24'b000000000000000000000001, 
24'b000000001100000000100101, 
24'b000000000000000000000000, 
24'b000000001101000000100101, 
24'b000000000000000000000000, 
24'b000000001101000000100100, 
24'b000000000000000000000001, 
24'b000000001011000000100011, 
24'b000000000000000000000000, 
24'b000000001100000000100011, 
24'b000000000000000000000000, 
24'b000000001100000000100010, 
24'b000000000000000000000000, 
24'b000000001100000000100001, 
24'b000000000000000000000001, 
24'b000000001011000000100001, 
24'b000000000000000000000000, 
24'b000000001011000000100000, 
24'b000000000000000000000000, 
24'b000000001011000000100000, 
24'b000000000000000000000000, 
24'b000000001010000000011111, 
24'b000000000000000000000000, 
24'b000000001010000000011111, 
24'b000000000000000000000000, 
24'b000000001010000000011111, 
24'b000000000000000000000000, 
24'b000000001010000000011110, 
24'b000000000000000000000000, 
24'b000000001010000000011101, 
24'b000000000000000000000000, 
24'b000000001010000000011101, 
24'b111111111111000000000000, 
24'b000000001010000000011100, 
24'b000000000000000000000000, 
24'b000000001010000000011100, 
24'b111111111111000000000000, 
24'b000000001001000000011011, 
24'b000000000000000000000000, 
24'b000000001001000000011011, 
24'b000000000001111111111111, 
24'b000000001010000000011011, 
24'b000000000000000000000000, 
24'b000000001001000000011011, 
24'b000000000000000000000000, 
24'b000000001001000000011010, 
24'b000000000000000000000000, 
24'b000000001001000000011010, 
24'b000000000000000000000000, 
24'b000000001010000000011001, 
24'b000000000000000000000000, 
24'b000000001001000000011001, 
24'b000000000000000000000000, 
24'b000000001001000000011001, 
24'b000000000000000000000000, 
24'b000000001001000000011000, 
24'b000000000000000000000000, 
24'b000000001001000000011000, 
24'b000000000000000000000000, 
24'b000000001000000000010111, 
24'b000000000000000000000000, 
24'b000000001000000000011000, 
24'b000000000000000000000000, 
24'b000000001000000000010111, 
24'b000000000000111111111111, 
24'b000000001001000000010111, 
24'b000000000000000000000000, 
24'b000000001000000000010110, 
24'b000000000000000000000000, 
24'b000000001000000000010110, 
24'b000000000000000000000000, 
24'b000000001001000000010110, 
24'b000000000000000000000000, 
24'b000000001000000000010110, 
24'b000000000000000000000000, 
24'b000000001000000000010110, 
24'b000000000000000000000000, 
24'b000000000111000000010110, 
24'b000000000000111111111111, 
24'b000000001000000000010101, 
24'b000000000000111111111111, 
24'b000000001001000000010101, 
24'b000000000000000000000000, 
24'b000000001000000000010101, 
24'b000000000000000000000000, 
24'b000000001000000000010101, 
24'b000000000000111111111111, 
24'b000000001000000000010100, 
24'b000000000000000000000000, 
24'b000000001000000000010100, 
24'b000000000000000000000000, 
24'b000000001000000000010011, 
24'b000000000001000000000000, 
24'b000000001000000000010101, 
24'b111111111111000000000000, 
24'b000000001000000000010011, 
24'b111111111111000000000000, 
24'b000000000111000000010010, 
24'b000000000001000000000000, 
24'b000000001000000000010011, 
24'b000000000000000000000001, 
24'b000000000111000000010010, 
24'b000000000000111111111111, 
24'b000000001000000000010011, 
24'b000000000000000000000000, 
24'b000000001000000000010010, 
24'b000000000000000000000000, 
24'b000000000111000000010010, 
24'b000000000000111111111111, 
24'b000000001000000000010010, 
24'b000000000001111111111111, 
24'b000000001001000000010010, 
24'b000000000000000000000000, 
24'b000000001001000000010010, 
24'b000000000000000000000001, 
24'b000000001000000000010010, 
24'b000000000001000000000000, 
24'b000000001000000000010010, 
24'b111111111111000000000000, 
24'b000000000111000000010001, 
24'b000000000001000000000000, 
24'b000000001000000000010010, 
24'b000000000000000000000000, 
24'b000000000111000000010001, 
24'b000000000000000000000000, 
24'b000000001000000000010001, 
24'b000000000000000000000000, 
24'b000000001000000000010001, 
24'b000000000000000000000000, 
24'b000000000111000000010001, 
24'b000000000000000000000000, 
24'b000000000111000000010001, 
24'b000000000000000000000000, 
24'b000000001000000000010000, 
24'b000000000000111111111111, 
24'b000000001000000000010001, 
24'b000000000000000000000000, 
24'b000000000111000000010000, 
24'b000000000000111111111111, 
24'b000000001001000000010000, 
24'b000000000000000000000000, 
24'b000000001000000000010000, 
24'b111111111111000000000001, 
24'b000000001000000000010000, 
24'b000000000000000000000000, 
24'b000000001000000000001111, 
24'b000000000000000000000000, 
24'b000000001000000000001111, 
24'b000000000000000000000001, 
24'b000000000111000000001111, 
24'b000000000000000000000000, 
24'b000000000111000000001111, 
24'b000000000000111111111111, 
24'b000000001001000000001111, 
24'b000000000000000000000001, 
24'b000000000111000000001111, 
24'b000000000000000000000001, 
24'b000000000111000000001110, 
24'b000000000001000000000000, 
24'b000000001000000000001111, 
24'b000000000001000000000000, 
24'b000000001000000000001111, 
24'b000000000000000000000001, 
24'b000000000111000000001111, 
24'b000000000000000000000001, 
24'b000000000111000000001110, 
24'b000000000000000000000000, 
24'b000000001000000000001110, 
24'b000000000000000000000001, 
24'b000000000111000000001111, 
24'b111111111111000000000000, 
24'b000000000111000000001110, 
24'b000000000001000000000000, 
24'b000000000111000000001111, 
24'b111111111111000000000000, 
24'b000000000111000000001101, 
24'b000000000001111111111111, 
24'b000000000111000000001110, 
24'b000000000000111111111111, 
24'b000000001000000000001110, 
24'b000000000000000000000000, 
24'b000000001000000000001101, 
24'b000000000000000000000000, 
24'b000000001000000000001110, 
24'b000000000000000000000000, 
24'b000000000111000000001110, 
24'b111111111111000000000000, 
24'b000000001000000000001101, 
24'b000000000000000000000000, 
24'b000000001000000000001101, 
24'b000000000000000000000000, 
24'b000000000111000000001101, 
24'b000000000000000000000000, 
24'b000000000111000000001101, 
24'b000000000000000000000000, 
24'b000000001000000000001101, 
24'b000000000000000000000000, 
24'b000000000111000000001101, 
24'b000000000000000000000000, 
24'b000000001000000000001100, 
24'b000000000000000000000000, 
24'b000000001000000000001100, 
24'b000000000000000000000000, 
24'b000000000111000000001101, 
24'b000000000000000000000000, 
24'b000000000111000000001100, 
24'b000000000000111111111111, 
24'b000000001000000000001100, 
24'b000000000000000000000000, 
24'b000000001000000000001100, 
24'b000000000000000000000000, 
24'b000000000111000000001100, 
24'b000000000000000000000000, 
24'b000000000111000000001100, 
24'b000000000000000000000000, 
24'b000000000111000000001100, 
24'b000000000000000000000000, 
24'b000000000111000000001100, 
24'b000000000000000000000000, 
24'b000000000111000000001100, 
24'b000000000000000000000000, 
24'b000000001000000000001011, 
24'b000000000001000000000000, 
24'b000000001000000000001101, 
24'b000000000000000000000000, 
24'b000000001000000000001100, 
24'b111111111111000000000001, 
24'b000000000111000000001011, 
24'b000000000000000000000000, 
24'b000000000111000000001011, 
24'b000000000000000000000000, 
24'b000000000110000000001100, 
24'b000000000000111111111111, 
24'b000000000111000000001011, 
24'b000000000001111111111111, 
24'b000000001000000000001100, 
24'b000000000000000000000000, 
24'b000000001000000000001011, 
24'b000000000000000000000001, 
24'b000000000111000000001011, 
24'b000000000000111111111111, 
24'b000000001000000000001011, 
24'b000000000001000000000000, 
24'b000000001000000000001011, 
24'b000000000000000000000000, 
24'b000000001000000000001011, 
24'b000000000000000000000000, 
24'b000000001000000000001011, 
24'b000000000000000000000000, 
24'b000000001000000000001011, 
24'b000000000000000000000000, 
24'b000000001000000000001011, 
24'b000000000000000000000000, 
24'b000000001000000000001011, 
24'b000000000000000000000000, 
24'b000000000111000000001010, 
24'b000000000001111111111111, 
24'b000000001000000000001011, 
24'b000000000001000000000000, 
24'b000000001000000000001011, 
24'b000000000000111111111111, 
24'b000000001000000000001011, 
24'b000000000000111111111111, 
24'b000000001001000000001011, 
24'b000000000000000000000001, 
24'b000000001000000000001011, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b000000000001000000000000, 
24'b000000001001000000001011, 
24'b111111111111000000000001, 
24'b000000000111000000001010, 
24'b000000000000111111111111, 
24'b000000001001000000001010, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b111111111111000000000000, 
24'b000000001000000000001010, 
24'b000000000000000000000000, 
24'b000000001000000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b000000000001000000000000, 
24'b000000001000000000001010, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b000000000000000000000000, 
24'b000000001000000000001001, 
24'b000000000001000000000000, 
24'b000000001000000000001010, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b000000000000111111111111, 
24'b000000001000000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001010, 
24'b000000000000000000000001, 
24'b000000000111000000001010, 
24'b000000000000111111111111, 
24'b000000001000000000001010, 
24'b111111111111000000000000, 
24'b000000001001000000001001, 
24'b000000000000000000000001, 
24'b000000001000000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001001, 
24'b000000000000111111111111, 
24'b000000001001000000001001, 
24'b000000000000000000000000, 
24'b000000001001000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001000, 
24'b000000000000000000000000, 
24'b000000001000000000001000, 
24'b000000000000000000000000, 
24'b000000001001000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001000, 
24'b000000000000111111111111, 
24'b000000001001000000001000, 
24'b000000000000000000000000, 
24'b000000001001000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001000, 
24'b000000000001000000000000, 
24'b000000001000000000001001, 
24'b000000000000111111111111, 
24'b000000001001000000001000, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000001000000000000, 
24'b000000001001000000001001, 
24'b000000000000000000000000, 
24'b000000001001000000001000, 
24'b000000000000000000000000, 
24'b000000001001000000001000, 
24'b000000000000000000000000, 
24'b000000001001000000001001, 
24'b000000000000000000000001, 
24'b000000001000000000001001, 
24'b111111111111000000000000, 
24'b000000001000000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000001000, 
24'b000000000001000000000000, 
24'b000000001000000000001001, 
24'b000000000000000000000000, 
24'b000000001000000000001000, 
24'b000000000000111111111111, 
24'b000000001010000000001000, 
24'b000000000000000000000001, 
24'b000000001001000000001000, 
24'b000000000000000000000001, 
24'b000000001000000000001000, 
24'b111111111111000000000000, 
24'b000000001000000000000111, 
24'b000000000000111111111111, 
24'b000000001001000000000111, 
24'b000000000000111111111111, 
24'b000000001001000000000111, 
24'b000000000001000000000000, 
24'b000000001001000000001001, 
24'b111111111111000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001000000000001000, 
24'b000000000000111111111111, 
24'b000000001010000000000111, 
24'b000000000000000000000001, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001000000000000111, 
24'b000000000000111111111111, 
24'b000000001001000000000111, 
24'b000000000001000000000000, 
24'b000000001010000000001000, 
24'b111111111111000000000001, 
24'b000000001001000000000111, 
24'b000000000000000000000001, 
24'b000000001000000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000001, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b111111111111000000000000, 
24'b000000001000000000000110, 
24'b000000000000111111111111, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000111111111111, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000111111111111, 
24'b000000001001000000000111, 
24'b000000000000111111111111, 
24'b000000001010000000000111, 
24'b111111111111000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000111, 
24'b000000000000000000000001, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000111111111111, 
24'b000000001010000000000101, 
24'b000000000000000000000001, 
24'b000000001001000000000110, 
24'b000000000000111111111111, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000001000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000111111111111, 
24'b000000001010000000000101, 
24'b000000000001000000000000, 
24'b000000001010000000000110, 
24'b000000000001111111111111, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000001000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b0_00000001010000000000110,
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000111111111111, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b111111111111000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000100111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000100111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000001, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101000000000000, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000111111111111, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000111111111111, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000101111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000001, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000111111111111, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000001000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000111111111111, 
24'b000000001000111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000001000111111111110, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000001000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000001000000000000, 
24'b000000001000111111111110, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111100, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001000111111111101, 
24'b000000000000111111111111, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111101, 
24'b000000000001000000000000, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000001000000000000, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111101, 
24'b111111111111000000000000, 
24'b000000001001111111111101, 
24'b111111111111000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000001, 
24'b000000001001111111111101, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000001, 
24'b000000001010111111111100, 
24'b000000000000000000000001, 
24'b000000001001111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001010111111111011, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001011111111111100, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001010111111111100, 
24'b000000000000000000000000, 
24'b000000001010111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111100, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111011, 
24'b000000000000000000000000, 
24'b000000001100111111111011, 
24'b000000000000000000000000, 
24'b000000001100111111111011, 
24'b000000000000000000000000, 
24'b000000001100111111111011, 
24'b000000000000000000000000, 
24'b000000001100111111111011, 
24'b000000000000000000000000, 
24'b000000001100111111111011, 
24'b000000000000000000000000, 
24'b000000001011111111111010, 
24'b000000000000000000000000, 
24'b000000001100111111111011, 
24'b000000000000000000000000, 
24'b000000001100111111111010, 
24'b000000000000000000000000, 
24'b000000001100111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001100111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001110111111111010, 
24'b000000000000000000000000, 
24'b000000001101111111111010, 
24'b000000000000000000000000, 
24'b000000001110111111111010, 
24'b000000000000000000000000, 
24'b000000001110111111111010, 
24'b000000000000000000000000, 
24'b000000001110111111111010, 
24'b000000000000000000000000, 
24'b000000001110111111111001, 
24'b000000000000000000000001, 
24'b000000001101111111111001, 
24'b000000000000000000000000, 
24'b000000001110111111111001, 
24'b000000000001000000000000, 
24'b000000001110111111111010, 
24'b000000000001000000000000, 
24'b000000001110111111111010, 
24'b000000000000000000000000, 
24'b000000001110111111111010, 
24'b000000000000000000000000, 
24'b000000001111111111111001, 
24'b000000000000000000000000, 
24'b000000001111111111111010, 
24'b000000000000000000000000, 
24'b000000001111111111111010, 
24'b000000000000000000000000, 
24'b000000001111111111111001, 
24'b000000000000000000000000, 
24'b000000001111111111111001, 
24'b000000000000000000000000, 
24'b000000001111111111111001, 
24'b000000000000000000000000, 
24'b000000010000111111111001, 
24'b000000000000000000000000, 
24'b000000010000111111111001, 
24'b000000000000000000000000, 
24'b000000010000111111111001, 
24'b000000000000000000000000, 
24'b000000010000111111111001, 
24'b111111111111000000000000, 
24'b000000010000111111111000, 
24'b000000000000000000000000, 
24'b000000010001111111111000, 
24'b000000000000000000000000, 
24'b000000010001111111111000, 
24'b000000000000000000000000, 
24'b000000010001111111111000, 
24'b000000000000000000000000, 
24'b000000010001111111111000, 
24'b000000000000000000000000, 
24'b000000010001111111111000, 
24'b000000000000000000000000, 
24'b000000010010111111111000, 
24'b000000000000000000000000, 
24'b000000010010111111111000, 
24'b000000000000000000000000, 
24'b000000010010111111111000, 
24'b111111111111000000000000, 
24'b000000010010111111110111, 
24'b000000000000000000000000, 
24'b000000010011111111110111, 
24'b000000000000000000000001, 
24'b000000010010111111110111, 
24'b000000000000000000000000, 
24'b000000010011111111110111, 
24'b000000000001000000000000, 
24'b000000010011111111111000, 
24'b000000000000000000000000, 
24'b000000010011111111110111, 
24'b000000000000111111111111, 
24'b000000010100111111110111, 
24'b000000000000000000000000, 
24'b000000010100111111110111, 
24'b000000000000000000000000, 
24'b000000010101111111110111, 
24'b000000000000000000000000, 
24'b000000010100111111110111, 
24'b000000000000000000000000, 
24'b000000010101111111110111, 
24'b000000000000000000000000, 
24'b000000010101111111110111, 
24'b000000000000000000000000, 
24'b000000010110111111110111, 
24'b000000000000000000000000, 
24'b000000010110111111110110, 
24'b000000000000000000000001, 
24'b000000010110111111110110, 
24'b000000000000000000000000, 
24'b000000010111111111110110, 
24'b000000000000000000000000, 
24'b000000010111111111110110, 
24'b000000000000000000000000, 
24'b000000011000111111110110, 
24'b000000000000000000000000, 
24'b000000011000111111110110, 
24'b000000000000000000000000, 
24'b000000011001111111110101, 
24'b000000000000000000000000, 
24'b000000011001111111110110, 
24'b000000000000000000000000, 
24'b000000011001111111110110, 
24'b000000000000000000000000, 
24'b000000011010111111110101, 
24'b000000000000000000000000, 
24'b000000011011111111110110, 
24'b000000000000000000000000, 
24'b000000011011111111110101, 
24'b000000000000000000000000, 
24'b000000011100111111110101, 
24'b000000000000000000000000, 
24'b000000011100111111110101, 
24'b000000000000000000000000, 
24'b000000011101111111110101, 
24'b000000000000000000000000, 
24'b000000011110111111110101, 
24'b000000000000000000000000, 
24'b000000011110111111110100, 
24'b000000000000111111111111, 
24'b000000011111111111110100, 
24'b000000000000000000000000, 
24'b000000100000111111110100, 
24'b000000000000000000000001, 
24'b000000100000111111110100, 
24'b000000000000000000000000, 
24'b000000100001111111110100, 
24'b000000000000000000000000, 
24'b000000100010111111110011, 
24'b000000000000000000000000, 
24'b000000100011111111110011, 
24'b000000000000000000000000, 
24'b000000100100111111110011, 
24'b000000000000000000000000, 
24'b000000100101111111110011, 
24'b000000000000000000000000, 
24'b000000100110111111110011, 
24'b000000000000000000000000, 
24'b000000101000111111110011, 
24'b000000000000000000000000, 
24'b000000101001111111110011, 
24'b000000000000000000000000, 
24'b000000101010111111110010, 
24'b000000000001000000000000, 
24'b000000101100111111110011, 
24'b000000000000000000000000, 
24'b000000101110111111110010, 
24'b000000000000000000000001, 
24'b000000101110111111110001, 
24'b000000000000111111111111, 
24'b000000110001111111110001, 
24'b000000000000000000000000, 
24'b000000110010111111110001, 
24'b000000000000000000000000, 
24'b000000110101111111110000, 
24'b000000000000000000000000, 
24'b000000110111111111110000, 
24'b000000000000000000000000, 
24'b000000111001111111101111, 
24'b000000000000000000000000, 
24'b000000111101111111101111, 
24'b000000000000000000000000, 
24'b000000111111111111101110, 
24'b000000000001111111111111, 
24'b000001000011111111101110, 
24'b000000000000000000000000, 
24'b000001000110111111101100, 
24'b000000000000111111111111, 
24'b000001001011111111101011, 
24'b000000000000000000000000, 
24'b000001010000111111101010, 
24'b000000000000000000000000, 
24'b000001010101111111101000, 
24'b000000000000000000000000, 
24'b000001011011111111100101, 
24'b000000000000000000000000, 
24'b000001100010111111100010, 
24'b000000000000000000000000, 
24'b000001101010111111011101, 
24'b000000000000000000000000, 
24'b000001110100111111010110, 
24'b000000000000000000000000, 
24'b000001111110111111001100, 
24'b000000000000000000000000, 
24'b000010001011111110111010, 
24'b000000000000000000000000, 
24'b000010010110111110011011, 
24'b000000000000000000000000, 
24'b000010010100111101010000, 
24'b000000000000000000000000, 
24'b111111010001110111110101, 
24'b001011010110110100101011, 
24'b010100000101000010010000, 
24'b001011010101001011010110, 
24'b000110110011010000000111, 
24'b110100101011001011010110, 
24'b000001000001110111111110, 
24'b001011010110001011010101, 
24'b110100111111001110001011, 
24'b110100101011110100101011, 
24'b001111111011110111011011, 
24'b001011010101001011010101, 
24'b000100100010001110010100, 
24'b110100101011001011010110, 
24'b000000110001111000010000, 
24'b001011010101001011010110, 
24'b111101110001010000100001, 
24'b110100101011001011010110, 
24'b111001111100000010100001, 
24'b110100101010001011010110, 
24'b101110010111110100111011, 
24'b001011010110110100101011, 
24'b001000111010001111000010, 
24'b110100101010001011010101, 
24'b111011101110000010110110, 
24'b110100101010001011010101, 
24'b101110001111111101111110, 
24'b110100101010110100101011, 
24'b000111101000111000101100, 
24'b110100101011001011010110, 
24'b111001001011101010101100, 
24'b001011010110001011010110, 
24'b101001001100111010100010, 
24'b001011010101110100101011, 
24'b110111100111000010101110, 
24'b001011010101110100101010, 
24'b111101100000010010100001, 
24'b110100101011110100101011, 
24'b000011010001000100011100, 
24'b110100101010110100101011, 
24'b010001010110111111000011, 
24'b110100101010001011010110, 
24'b000000100110111001111111, 
24'b110100101010001011010101, 
24'b110000001101101101011111, 
24'b001011010101110100101011, 
24'b111111111011000111000101, 
24'b110100101011110100101011, 
24'b001111001010111000100110, 
24'b110100101010001011010101, 
24'b111000001000101000011111, 
24'b001011010110110100101010, 
24'b010000011001110110101110, 
24'b001011010101001011010110, 
24'b000011011011111100010011, 
24'b001011010101001011010101, 
24'b111110000111000001100100, 
24'b001011010101001011010110, 
24'b111000011111001110011000, 
24'b110100101011001011010110, 
24'b101010001011110101101110, 
24'b001011010110110100101010, 
24'b111001101011001011100101, 
24'b110100101010110100101010, 
24'b000001011001110100011110, 
24'b001011010110110100101010, 
24'b010000011010001010111010, 
24'b110100101010001011010110, 
24'b000000011011110100001000, 
24'b001011010110001011010101, 
24'b110001011101001010110110, 
24'b110100101010110100101011, 
24'b001001010100110100011101, 
24'b001011010110001011010101, 
24'b110011001010001100001111, 
24'b110100101011110100101011, 
24'b001010010010111101011110, 
24'b110100101010001011010101, 
24'b110100010001101110100101, 
24'b001011010101110100101011, 
24'b001100100100000101111001, 
24'b110100101010001011010110, 
24'b111110111111101110000110, 
24'b001011010101001011010110, 
24'b110111110100111100011100, 
24'b001011010101001011010110, 
24'b101000100101001010011000, 
24'b110100101011110100101010, 
24'b110111000100110000111011, 
24'b001011010110110100101011, 
24'b111100110010111110110000, 
24'b001011010101110100101010, 
24'b000010010100001100110000, 
24'b110100101010110100101011, 
24'b010000000001110100001111, 
24'b001011010110001011010101, 
24'b111110101110001001110001, 
24'b110100101011001011010110, 
24'b101101011101110001011101, 
24'b001011010101110100101010, 
24'b111011010101111111111101, 
24'b001011010101110100101011, 
24'b000001100110001111010011, 
24'b110100101010110100101011, 
24'b001110010101111110111010, 
24'b110100101011001011010101, 
24'b110100101001101111001101, 
24'b001011010101110100101011, 
24'b000010101111000101110011, 
24'b110100101011110100101011, 
24'b010010000001101101000110, 
24'b001011010101001011010110, 
24'b000001110001111001100010, 
24'b001011010110001011010101, 
24'b110010011000111110001001, 
24'b001011010101110100101011, 
24'b001001100010000010100011, 
24'b001011010101001011010110, 
24'b110001110111001110010100, 
24'b110100101011110100101010, 
24'b000000101110110011101001, 
24'b001011010110110100101010, 
24'b010000001110111111111101, 
24'b001011010101001011010101, 
24'b111111101111000110001000, 
24'b001011010101001011010101, 
24'b101111000101010100010110, 
24'b110100101010110100101011, 
24'b111101100111000100100010, 
24'b110100101010110100101011, 
24'b000100111100111100010101, 
24'b110100101011110100101010, 
24'b010100000100101100100000, 
24'b001011010101001011010110, 
24'b000101010010111010100110, 
24'b001011010101001011010101, 
24'b111111000011000000000111, 
24'b001011010101001011010101, 
24'b111000101110000101100011, 
24'b001011010110001011010110, 
24'b101001100011010011010111, 
24'b110100101011110100101011, 
24'b110111110100000010100010, 
24'b110100101010110100101011, 
24'b111100111100110010101111, 
24'b001011010101110100101011, 
24'b000000110101001001100011, 
24'b110100101011110100101011, 
24'b000101011000110001011111, 
24'b001011010101110100101010, 
24'b010001101110111111101010, 
24'b001011010101001011010110, 
24'b111000101000001101100011, 
24'b110100101011110100101011, 
24'b001101110100110100001011, 
24'b001011010110001011010101, 
24'b110101001001000010010100, 
24'b001011010101110100101010, 
24'b000010100100010001011010, 
24'b110100101011110100101011, 
24'b001001101101000000101101, 
24'b110100101010110100101011, 
24'b011001000101101111111111, 
24'b001011010110001011010110, 
24'b001010111110111111000110, 
24'b001011010101001011010110, 
24'b000110000100001101001110, 
24'b110100101010001011010101, 
24'b000010101001110011110100, 
24'b001011010101001011010101, 
24'b111111010111000001100110, 
24'b001011010101001011010110, 
24'b111010111100001111011101, 
24'b110100101011001011010101, 
24'b101101111010110110010000, 
24'b001011010101110100101011, 
24'b111111101110000100110010, 
24'b001011010110110100101011, 
24'b010001100010010100101111, 
24'b110100101010001011010101, 
24'b000100100001000110000001, 
24'b110100101011001011010110, 
24'b000000000110111111001001, 
24'b110100101010001011010101, 
24'b111100110101110001111000, 
24'b001011010110001011010101, 
24'b111001011100001011000100, 
24'b110100101011001011010110, 
24'b110100101000111100011001, 
24'b110100101010001011010101, 
24'b100110110010101100010101, 
24'b001011010101110100101010, 
24'b110111001000111010111101, 
24'b001011010101110100101010, 
24'b000101101110000010000000, 
24'b001011010110001011010101, 
24'b101100001100010000010100, 
24'b110100101011110100101011, 
24'b111000110001111111011001, 
24'b110100101011110100101010, 
24'b111110011001101110100100, 
24'b001011010101110100101011, 
24'b001010011100111101100000, 
24'b001011010110001011010101, 
24'b101111100101001011011000, 
24'b110100101010110100101011, 
24'b111011000110110001011101, 
24'b001011010110110100101010, 
24'b111111000001111101111110, 
24'b001011010110110100101011, 
24'b000010001111000011110101, 
24'b001011010101110100101011, 
24'b000110011001010000100110, 
24'b110100101011110100101010, 
24'b010010100100110111110000, 
24'b001011010110001011010110, 
24'b111001011110001101010101, 
24'b110100101011110100101010, 
24'b001111000011110101111010, 
24'b001011010101001011010110, 
24'b110111110001001011111000, 
24'b110100101011110100101011, 
24'b001110001000110100011011, 
24'b001011010110001011010110, 
24'b110111011110001001111110, 
24'b110100101010110100101011, 
24'b001110111011110001000000, 
24'b001011010101001011010110, 
24'b111111101001111101100001, 
24'b001011010101001011010101, 
24'b101111010111000010011011, 
24'b001011010110110100101010, 
24'b111110000100000111100110, 
24'b001011010101110100101010, 
24'b000101011010010101001101, 
24'b110100101011110100101010, 
24'b010100011010000100000111, 
24'b110100101011001011010110, 
24'b000101010000110011100000, 
24'b001011010110001011010101, 
24'b111101101111000011010000, 
24'b001011010101001011010110, 
24'b101110110101010011010101, 
24'b110100101011110100101010, 
24'b111110110101000100010011, 
24'b110100101011110100101010, 
24'b001101101001111100011101, 
24'b110100101010001011010101, 
24'b110100111101101100110000, 
24'b001011010110110100101010, 
24'b000011110110111010110001, 
24'b001011010110110100101011, 
24'b010100000000111111110110, 
24'b001011010110001011010101, 
24'b000101011101000011110101, 
24'b001011010101001011010101, 
24'b111110101000001000101100, 
24'b001011010110001011010110, 
24'b110001001110010110001011, 
24'b110100101011110100101011, 
24'b001001100100000100111001, 
24'b110100101011001011010110, 
24'b110011100001110011110110, 
24'b001011010101110100101011, 
24'b001010011110000010001100, 
24'b001011010101001011010101, 
24'b110011111010001001011000, 
24'b001011010110110100101011, 
24'b001010100101011000010011, 
24'b110100101010001011010110, 
24'b110011110001001000100111, 
24'b110100101011110100101010, 
24'b001010000011111010011111, 
24'b001011010110001011010101, 
24'b110010001111010100100001, 
24'b110100101010110100101011, 
24'b000001000100001000101011, 
24'b110100101011110100101011, 
24'b010000101000000100101111, 
24'b110100101010001011010101, 
24'b000000010100000001110111, 
24'b110100101010001011010101, 
24'b110000000000111110111111, 
24'b110100101011110100101010, 
24'b111111100111111011000101, 
24'b110100101010110100101011, 
24'b001110100010101111010010, 
24'b001011010101001011010101, 
24'b110110111110001001011010, 
24'b110100101011110100101011, 
24'b001110001101111011011011, 
24'b110100101010001011010101, 
24'b111110111001101011111000, 
24'b001011010101001011010101, 
24'b101110110000111010111101, 
24'b001011010101110100101010, 
24'b111110001010000010010010, 
24'b001011010110110100101011, 
24'b001100011110010000010101, 
24'b110100101010001011010101, 
24'b110011001010111000111011, 
24'b001011010101110100101011, 
24'b000000111111010000111110, 
24'b110100101011110100101010, 
24'b001110110001000011110000, 
24'b110100101010001011010101, 
24'b110101010101111101100101, 
24'b110100101011110100101011, 
24'b000011010001110000110111, 
24'b001011010110110100101011, 
24'b010001100000001010101010, 
24'b110100101011001011010110, 
24'b111001001101111101000010, 
24'b110100101011110100101011, 
24'b001100100000110001101110, 
24'b000000000000000000000000, 
24'b001101111001110001100110, 
24'b001011010110001011010101, 
24'b000011110000111100010000, 
24'b001011010101001011010110, 
24'b111101010000000011000011, 
24'b001011010110001011010110, 
24'b101110110010010001111010, 
24'b110100101011110100101011, 
24'b111110111111000010101110, 
24'b110100101010110100101010, 
24'b001101111001111011010101, 
24'b110100101010001011010101, 
24'b110101001110101101001100, 
24'b001011010101110100101010, 
24'b000011111101000100011000, 
24'b110100101010110100101011, 
24'b010011101011101011111000, 
24'b001011010110001011010101, 
24'b000011101100111000010101, 
24'b001011010110001011010101, 
24'b110011111010111100100110, 
24'b001011010101110100101011, 
24'b000100011100111111110110, 
24'b001011010110110100101010, 
24'b010101011110000011101101, 
24'b001011010110001011010110, 
24'b000111110000001111000100, 
24'b110100101011001011010110, 
24'b000010011011110011111100, 
24'b001011010101001011010101, 
24'b111101001001111111011100, 
24'b001011010110001011010101, 
24'b101111100011000011101101, 
24'b001011010110110100101011, 
24'b000000110101001000001101, 
24'b001011010110110100101010, 
24'b010001110110010100100010, 
24'b110100101010001011010101, 
24'b000010110111111011100100, 
24'b001011010110001011010101, 
24'b110100101011010001001110, 
24'b110100101010110100101011, 
24'b001101010011111010000010, 
24'b001011010101001011010101, 
24'b111000001110010000011101, 
24'b110100101011110100101010, 
24'b010001011100111001110010, 
24'b001011010110001011010101, 
24'b000101000001010000101101, 
24'b110100101011001011010110, 
24'b111111100111111010101110, 
24'b001011010101001011010110, 
24'b110011110000010011001110, 
24'b110100101010110100101011, 
24'b001110110010000110001001, 
24'b110100101011001011010110, 
24'b000011011010111111111111, 
24'b110100101010001011010110, 
24'b111111100100110011000011, 
24'b001011010110001011010110, 
24'b111100010010001011111001, 
24'b110100101011001011010101, 
24'b110111111000110110100111, 
24'b001011010110001011010101, 
24'b101010101010001111001100, 
24'b110100101010110100101010, 
24'b111011111010000001001110, 
24'b110100101010110100101011, 
24'b001100000010110011011010, 
24'b001011010101001011010110, 
24'b110101100100001100110110, 
24'b110100101011110100101011, 
24'b001110001000111110111010, 
24'b110100101011001011010101, 
24'b000001001101110000101000, 
24'b001011010101001011010110, 
24'b111011001000001000101000, 
24'b110100101010001011010101, 
24'b101110001110110010001011, 
24'b001011010110110100101011, 
24'b000110111011001000011000, 
24'b110100101010001011010110, 
24'b110001001010101111111100, 
24'b001011010110110100101011, 
24'b001000010110111100110111, 
24'b001011010110001011010110, 
24'b110001111101000010000111, 
24'b001011010101110100101010, 
24'b001000101010000111011101, 
24'b001011010101001011010110, 
24'b110001010001010100101101, 
24'b110100101011110100101011, 
24'b000000101011111101000001, 
24'b001011010101110100101011, 
24'b010001001001010101001000, 
24'b110100101011001011010110, 
24'b000010110000001000011010, 
24'b110100101011001011010110, 
24'b111011110111000011111001, 
24'b110100101011001011010101, 
24'b101101101110000000011111, 
24'b110100101011110100101010, 
24'b111110110111111100111110, 
24'b110100101011110100101010, 
24'b010000001000111000000010, 
24'b110100101010001011010101, 
24'b000010011101101001111010, 
24'b001011010110001011010101, 
24'b111101000011111001010101, 
24'b001011010110001011010110, 
24'b110111100011000000100011, 
24'b001011010110001011010101, 
24'b101001100100001101111101, 
24'b110100101011110100101010, 
24'b111010001000110100110001, 
24'b001011010110110100101010, 
24'b001001011101000011010110, 
24'b001011010101001011010110, 
24'b110001110101010011000101, 
24'b110100101011110100101010, 
24'b001000001001000011011010, 
24'b110100101010001011010110, 
24'b110001000111110100110110, 
24'b001011010110110100101011, 
24'b000111001100001101111010, 
24'b110100101011001011010101, 
24'b101111000100111111101100, 
24'b110100101010110100101010, 
24'b111101010101110001001010, 
24'b001011010110110100101010, 
24'b001011011001001000110100, 
24'b110100101010001011010110, 
24'b110010001101110001010111, 
24'b001011010101110100101011, 
24'b000000100101000000000111, 
24'b001011010101110100101011, 
24'b001111111111001110100101, 
24'b110100101010001011010101, 
24'b111111110100110101110110, 
24'b001011010110001011010101, 
24'b110000011001000100110111, 
24'b001011010101110100101010, 
24'b000111011010010101010101, 
24'b110100101011001011010101, 
24'b101111010110000111011100, 
24'b110100101001110100101011, 
24'b111100110101000010001111, 
24'b110100101010110100101011, 
24'b000011101011111110000001, 
24'b110100101011110100101011, 
24'b010010001101111000101011, 
24'b110100101011001011010110, 
24'b000001111101101010010010, 
24'b001011010110001011010101, 
24'b110010111000111001010100, 
24'b001011010101110100101011, 
24'b001010110000111111100001, 
24'b001011010101001011010110, 
24'b110100111100000101100101, 
24'b001011010110110100101011, 
24'b001101010001010011111111, 
24'b110100101011001011010110, 
24'b111111101111000011110011, 
24'b110100101011001011010101, 
24'b111000101011110100110101, 
24'b001011010110001011010101, 
24'b101001101000001100110111, 
24'b110100101011110100101011, 
24'b111000011111110111001010, 
24'b001011010101110100101011, 
24'b111111010110001111100011, 
24'b110100101011110100101010, 
24'b001100101001000001100011, 
24'b110100101010001011010101, 
24'b110100000011110011110101, 
24'b001011010110110100101011, 
24'b001001100001001101101010, 
24'b110100101011001011010110, 
24'b110001001000000000111000, 
24'b110100101010110100101010, 
24'b111111011000111010011101, 
24'b110100101010110100101011, 
24'b001101101111101100010000, 
24'b001011010101001011010101, 
24'b110101110100111100111101, 
24'b001011010110110100101011, 
24'b001100110001001101001101, 
24'b110100101010001011010101, 
24'b111101001001111101000010, 
24'b110100101010001011010110, 
24'b101100100001101100011001, 
24'b001011010110110100101011, 
24'b111010101110111010101100, 
24'b001011010101110100101010, 
24'b000001010000000001010000, 
24'b001011010101110100101010, 
24'b001110011000001110010101, 
24'b110100101011001011010110, 
24'b110101101110110101011111, 
24'b001011010110110100101011, 
24'b001011010111001010101001, 
24'b110100101010001011010101, 
24'b110011111001110001100110, 
24'b001011010101110100101010, 
24'b001001100100111110000111, 
24'b001011010101001011010110, 
24'b110000111011000011000100, 
24'b001011010101110100101010, 
24'b111110001000001000001001, 
24'b001011010101110100101010, 
24'b000100110011010101000111, 
24'b110100101011110100101011, 
24'b010011010110111101000011, 
24'b001011010101001011010101, 
24'b000011110001010100011111, 
24'b110100101011001011010101, 
24'b111011110001000110000110, 
24'b110100101010001011010110, 
24'b101100001001111000010101, 
24'b001011010110110100101011, 
24'b111010100011010010011011, 
24'b110100101011110100101010, 
24'b000000111111000110011011, 
24'b110100101010110100101011, 
24'b001101100111000010000101, 
24'b110100101011001011010110, 
24'b110011011100111110010111, 
24'b110100101010110100101011, 
24'b000000000011111001011010, 
24'b110100101011110100101011, 
24'b000110011011101011011010, 
24'b001011010110110100101011, 
24'b010100101011111011000001, 
24'b001011010110001011010110, 
24'b000100010001000010100011, 
24'b001011010101001011010101, 
24'b110101001101010000100001, 
24'b110100101010110100101010, 
24'b001101110000111000101110, 
24'b001011010101001011010110, 
24'b111110110110001111011010, 
24'b110100101011001011010110, 
24'b101110111000111001010111, 
24'b001011010110110100101011, 
24'b111110011010010001101110, 
24'b110100101010110100101010, 
24'b001100110100000011110100, 
24'b110100101010001011010110, 
24'b110011101000110110010010, 
24'b001011010110110100101011, 
24'b000001100110010000010001, 
24'b110100101011110100101011, 
24'b001111101000000011001010, 
24'b110100101011001011010110, 
24'b110110100110110110010101, 
24'b001011010101110100101010, 
24'b000101010110010001001100, 
24'b110100101010110100101011, 
24'b010101100011000110000000, 
24'b110100101011001011010110, 
24'b000111010011000010101100, 
24'b110100101011001011010110, 
24'b000001100101000000100011, 
24'b110100101011001011010101, 
24'b111011111100111110101111, 
24'b110100101010001011010101, 
24'b101110000000111100111110, 
24'b110100101010110100101010, 
24'b111110111001111011000010, 
24'b110100101010110100101011, 
24'b001111011010111000100111, 
24'b110100101011001011010110, 
24'b111111110100110100110101, 
24'b110100101011001011010110, 
24'b110000101111101000101101, 
24'b001011010110110100101010, 
24'b000111111110000001011110, 
24'b110100101011001011010110, 
24'b101111111111101010101010, 
24'b001011010110110100101010, 
24'b111101011101111001110000, 
24'b001011010110110100101011, 
24'b000100000000001000100001, 
24'b110100101011110100101010, 
24'b010001011100110000011111, 
24'b001011010110001011010110, 
24'b111001010100000110001011, 
24'b110100101011110100101011, 
24'b001111110101101101101001, 
24'b001011010110001011010110, 
24'b111001110100111010111001, 
24'b001011010101110100101010, 
24'b010010100011000001011110, 
24'b001011010110001011010101, 
24'b000110000111001111101001, 
24'b110100101011001011010110, 
24'b000001101101111110110000, 
24'b110100101010001011010101, 
24'b111110010100101110000100, 
24'b001011010110001011010110, 
24'b111010101111111101010111, 
24'b001011010101001011010110, 
24'b110101101001001011111000, 
24'b110100101011001011010110, 
24'b100111001111110011100110, 
24'b001011010101110100101010, 
24'b110110000100001001001000, 
24'b110100101011110100101010, 
24'b111011110001110000100101, 
24'b001011010110110100101011, 
24'b000000100101111110001101, 
24'b001011010110110100101010, 
24'b001001011100001000011100, 
24'b000000000000000000000000, 
24'b000011011100000010111001, 
24'b000000000000000000000000, 
24'b000001111111000001101000, 
24'b000000000000000000000000, 
24'b000001010110000001000011, 
24'b000000000000000000000000, 
24'b000000111111000000101101, 
24'b000000000001000000000000, 
24'b000000110000000000100001, 
24'b000000000000000000000000, 
24'b000000100110000000011000, 
24'b000000000000000000000000, 
24'b000000100000000000010001, 
24'b000000000000000000000000, 
24'b000000011011000000001011, 
24'b000000000000000000000000, 
24'b000000010111000000001000, 
24'b000000000000000000000001, 
24'b000000010100000000000101, 
24'b000000000000000000000000, 
24'b000000010010000000000010, 
24'b000000000000000000000000, 
24'b000000010000000000000000, 
24'b111111111111000000000000, 
24'b000000001111111111111110, 
24'b000000000000000000000000, 
24'b000000001101111111111101, 
24'b000000000000000000000000, 
24'b000000001100111111111100, 
24'b000000000000111111111111, 
24'b000000001100111111111011, 
24'b000000000000000000000000, 
24'b000000001010111111111011, 
24'b000000000000000000000000, 
24'b000000001010111111111010, 
24'b000000000000000000000000, 
24'b000000001001111111111010, 
24'b000000000000000000000000, 
24'b000000001001111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000000111111111111001, 
24'b000000000000111111111111, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000000111111111111000, 
24'b000000000000000000000000, 
24'b000000000111111111111000, 
24'b000000000000000000000000, 
24'b000000000111111111111000, 
24'b000000000000000000000000, 
24'b000000000110111111111000, 
24'b000000000000000000000000, 
24'b000000000111111111111000, 
24'b000000000000000000000000, 
24'b000000000110111111111000, 
24'b000000000000000000000000, 
24'b000000000110111111111000, 
24'b000000000000000000000001, 
24'b000000000101111111111000, 
24'b000000000000000000000001, 
24'b000000000101111111111000, 
24'b000000000000000000000000, 
24'b000000000101111111111000, 
24'b000000000000000000000000, 
24'b000000000101111111111000, 
24'b000000000000000000000000, 
24'b000000000101111111111000, 
24'b000000000000000000000000, 
24'b000000000101111111111000, 
24'b000000000000000000000000, 
24'b000000000101111111111000, 
24'b000000000000000000000000, 
24'b000000000101111111111001, 
24'b000000000000000000000000, 
24'b000000000101111111111000, 
24'b000000000000000000000000, 
24'b000000000100111111111001, 
24'b000000000000000000000000, 
24'b000000000100111111111000, 
24'b000000000000000000000000, 
24'b000000000100111111111001, 
24'b000000000000000000000000, 
24'b000000000100111111111001, 
24'b000000000000000000000000, 
24'b000000000100111111111001, 
24'b000000000000000000000000, 
24'b000000000100111111111001, 
24'b000000000000000000000000, 
24'b000000000011111111111001, 
24'b000000000001000000000000, 
24'b000000000100111111111010, 
24'b000000000000000000000000, 
24'b000000000100111111111010, 
24'b000000000000000000000000, 
24'b000000000100111111111010, 
24'b000000000000000000000000, 
24'b000000000100111111111001, 
24'b000000000000000000000000, 
24'b000000000011111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111001, 
24'b000000000000000000000000, 
24'b000000000100111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b111111111111000000000000, 
24'b000000000011111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111010, 
24'b000000000000111111111111, 
24'b000000000100111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111010, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111011, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000010111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000010111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000010111111111100, 
24'b000000000000000000000000, 
24'b000000000010111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000011111111111100, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111100, 
24'b000000000000000000000000, 
24'b000000000010111111111100, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000011111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000011111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000011111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111100, 
24'b000000000001111111111111, 
24'b000000000011111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b111111111111000000000000, 
24'b000000000011111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000011111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000011111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000011111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111101, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000001000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b111111111111000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111110, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b111111111111000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b111111111111000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000111111111111, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000001, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000001000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010111111111111, 
24'b000000000001000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b111111111111000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000010000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000111111111111, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000111111111111, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000011111111111111, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000011000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b000000000100000000000000, 
24'b000000000000000000000000, 
24'b0_00000000100000000000000,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b111111111111000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b111111111111000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b111111111111000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000001, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000001000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000001, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000001, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111110, 
24'b111111111111000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000001000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000111111111111, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111101, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000001, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111101, 
24'b111111111111000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000001000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000001, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111100, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000001, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000110111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000111111111111, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000001000111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000001000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000001, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000001000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111011, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000001, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000001000111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111001, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000001000111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000001000111111111010, 
24'b000000000000000000000000, 
24'b000000000111111111111010, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111010, 
24'b111111111111000000000000, 
24'b000000000111111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000000111111111111001, 
24'b000000000000000000000000, 
24'b000000000111111111111001, 
24'b000000000000000000000000, 
24'b000000000111111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000000111111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b111111111111000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111001, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001000111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000001, 
24'b000000001001111111111000, 
24'b000000000000000000000001, 
24'b000000001000111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111111000, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001001111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b111111111111000000000000, 
24'b000000001010111111110110, 
24'b000000000000000000000000, 
24'b000000001010111111110110, 
24'b000000000000000000000000, 
24'b000000001010111111110110, 
24'b000000000000000000000000, 
24'b000000001010111111110111, 
24'b000000000000000000000000, 
24'b000000001010111111110110, 
24'b000000000000000000000000, 
24'b000000001010111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001011111111110110, 
24'b000000000000000000000000, 
24'b000000001100111111110101, 
24'b000000000000000000000000, 
24'b000000001011111111110101, 
24'b000000000000000000000000, 
24'b000000001011111111110101, 
24'b000000000000000000000000, 
24'b000000001011111111110101, 
24'b000000000000000000000000, 
24'b000000001100111111110101, 
24'b000000000000000000000000, 
24'b000000001100111111110101, 
24'b000000000000000000000000, 
24'b000000001100111111110101, 
24'b000000000000000000000000, 
24'b000000001100111111110101, 
24'b000000000000000000000000, 
24'b000000001100111111110101, 
24'b000000000000000000000000, 
24'b000000001101111111110101, 
24'b000000000000000000000000, 
24'b000000001101111111110101, 
24'b000000000000000000000000, 
24'b000000001100111111110101, 
24'b000000000000000000000000, 
24'b000000001101111111110101, 
24'b000000000000000000000000, 
24'b000000001101111111110101, 
24'b000000000000000000000000, 
24'b000000001101111111110101, 
24'b000000000000000000000000, 
24'b000000001101111111110100, 
24'b000000000000000000000000, 
24'b000000001101111111110100, 
24'b000000000000000000000000, 
24'b000000001101111111110100, 
24'b000000000000000000000000, 
24'b000000001101111111110101, 
24'b000000000000000000000000, 
24'b000000001110111111110100, 
24'b000000000000000000000000, 
24'b000000001110111111110100, 
24'b000000000000000000000000, 
24'b000000001110111111110100, 
24'b000000000000000000000000, 
24'b000000001110111111110100, 
24'b000000000000000000000000, 
24'b000000001110111111110100, 
24'b000000000000000000000000, 
24'b000000001111111111110011, 
24'b000000000000000000000000, 
24'b000000001111111111110100, 
24'b000000000000000000000000, 
24'b000000001111111111110011, 
24'b000000000000000000000000, 
24'b000000001111111111110011, 
24'b000000000000000000000000, 
24'b000000001111111111110011, 
24'b000000000000000000000000, 
24'b000000010000111111110011, 
24'b000000000000000000000000, 
24'b000000010000111111110011, 
24'b000000000000000000000000, 
24'b000000010000111111110011, 
24'b000000000000000000000000, 
24'b000000010000111111110011, 
24'b000000000000000000000000, 
24'b000000010000111111110011, 
24'b000000000000000000000000, 
24'b000000010001111111110011, 
24'b000000000000000000000000, 
24'b000000010001111111110011, 
24'b000000000000000000000000, 
24'b000000010001111111110011, 
24'b000000000000000000000000, 
24'b000000010001111111110010, 
24'b000000000000000000000000, 
24'b000000010010111111110010, 
24'b000000000000000000000000, 
24'b000000010010111111110011, 
24'b000000000000000000000000, 
24'b000000010011111111110010, 
24'b000000000000000000000000, 
24'b000000010011111111110010, 
24'b000000000000000000000000, 
24'b000000010011111111110010, 
24'b000000000000000000000000, 
24'b000000010011111111110010, 
24'b000000000000000000000000, 
24'b000000010100111111110010, 
24'b000000000000000000000000, 
24'b000000010100111111110001, 
24'b000000000000000000000000, 
24'b000000010101111111110001, 
24'b000000000000000000000000, 
24'b000000010101111111110010, 
24'b000000000000000000000000, 
24'b000000010110111111110001, 
24'b000000000000000000000000, 
24'b000000010110111111110001, 
24'b000000000000000000000000, 
24'b000000010110111111110001, 
24'b000000000000111111111111, 
24'b000000011000111111110001, 
24'b000000000000000000000000, 
24'b000000011000111111110001, 
24'b000000000000000000000000, 
24'b000000011000111111110000, 
24'b000000000000000000000000, 
24'b000000011001111111110000, 
24'b000000000000000000000000, 
24'b000000011010111111110000, 
24'b000000000000000000000000, 
24'b000000011010111111110000, 
24'b000000000000000000000000, 
24'b000000011011111111110000, 
24'b000000000000000000000000, 
24'b000000011100111111110000, 
24'b000000000000000000000000, 
24'b000000011101111111110000, 
24'b000000000000000000000000, 
24'b000000011101111111110000, 
24'b000000000000000000000000, 
24'b000000011111111111110000, 
24'b000000000000000000000000, 
24'b000000011111111111101111, 
24'b000000000000000000000000, 
24'b000000100000111111101111, 
24'b000000000000000000000000, 
24'b000000100001111111101111, 
24'b000000000000000000000000, 
24'b000000100010111111101111, 
24'b000000000000000000000001, 
24'b000000100011111111101111, 
24'b000000000000111111111111, 
24'b000000100101111111101111, 
24'b000000000000000000000000, 
24'b000000100110111111101110, 
24'b000000000000111111111111, 
24'b000000101000111111101101, 
24'b000000000000111111111111, 
24'b000000101010111111101101, 
24'b000000000000000000000000, 
24'b000000101011111111101101, 
24'b000000000000000000000000, 
24'b000000101101111111101101, 
24'b000000000000000000000000, 
24'b000000101111111111101100, 
24'b000000000000000000000000, 
24'b000000110010111111101100, 
24'b000000000000000000000000, 
24'b000000110100111111101011, 
24'b000000000000000000000000, 
24'b000000110111111111101011, 
24'b000000000000000000000000, 
24'b000000111001111111101010, 
24'b000000000000000000000000, 
24'b000000111101111111101010, 
24'b000000000000000000000000, 
24'b000001000000111111101001, 
24'b000000000000000000000000, 
24'b000001000101111111100111, 
24'b000000000000000000000000, 
24'b000001001001111111100101, 
24'b000000000000000000000000, 
24'b000001001111111111100100, 
24'b000000000000000000000000, 
24'b000001010101111111100001, 
24'b000000000000000000000000, 
24'b000001011011111111011110, 
24'b000000000000000000000000, 
24'b000001100100111111011001, 
24'b000000000000000000000000, 
24'b000001101101111111010010, 
24'b000000000000000000000000, 
24'b000001110111111111001000, 
24'b000000000000000000000000, 
24'b000010000011111110110111, 
24'b000000000000000000000000, 
24'b000010001110111110011000, 
24'b000000000000000000000000, 
24'b000010001100111101001110, 
24'b000000000000000000000000, 
24'b111111001011110111110110, 
24'b001011001111110100110001, 
24'b010011110011000010001011, 
24'b001011001111001011001111, 
24'b000110101001001111111010, 
24'b110100110001001011010000, 
24'b000000111001110111111110, 
24'b001011001111001011001111, 
24'b110100111110001101111110, 
24'b110100110001110100110001, 
24'b001111101011110111011100, 
24'b001011001111001011001111, 
24'b000100011000001110001000, 
24'b110100110001001011001111, 
24'b000000101010111000010001, 
24'b001011001111001011001111, 
24'b111101101011010000010100, 
24'b110100110001001011001111, 
24'b111001111001000010011100, 
24'b110100110000001011001111, 
24'b101110011011110100111110, 
24'b001011001111110100110001, 
24'b001000101110001110110101, 
24'b110100110000001011001111, 
24'b111011101010000010101111, 
24'b110100110001001011001111, 
24'b101110010001111101111011, 
24'b110100110001110100110001, 
24'b000111011101111000101101, 
24'b110100110001001011010000, 
24'b111001000111101010110100, 
24'b001011001111001011001111, 
24'b101001010001111010100001, 
24'b001011001111110100110001, 
24'b110111100100000010101000, 
24'b001011001111110100110000, 
24'b111101011001010010010011, 
24'b110100110001110100110000, 
24'b000011001001000100010101, 
24'b110100110001110100110010, 
24'b010001000101111110111111, 
24'b110100110001001011001111, 
24'b000000011101111001111110, 
24'b110100110001001011001111, 
24'b110000001110101101100110, 
24'b001011010000110100110001, 
24'b111111110011000110111110, 
24'b110100110001110100110001, 
24'b001110111001111000100110, 
24'b110100110001001011001111, 
24'b111000000100101000101000, 
24'b001011001111110100110001, 
24'b010000000111110110101111, 
24'b001011001111001011001111, 
24'b000011010000111100010001, 
24'b001011001111001011001111, 
24'b111101111111000001011111, 
24'b001011001111001011001111, 
24'b111000011011001110001100, 
24'b110100110001001011001111, 
24'b101010001111110101110000, 
24'b001011010000110100110001, 
24'b111001100111001011011010, 
24'b110100110001110100110001, 
24'b000001010000110100100001, 
24'b001011001111110100110001, 
24'b010000000111001010110000, 
24'b110100110001001011001111, 
24'b000000010001110100001011, 
24'b001011001111001011001111, 
24'b110001011100001010101100, 
24'b110100110001110100110000, 
24'b001001000101110100100000, 
24'b001011001111001011001111, 
24'b110011001000001100000101, 
24'b110100110001110100110001, 
24'b001010000011111101011100, 
24'b110100110001001011001111, 
24'b110100001111101110101011, 
24'b001011001111110100110001, 
24'b001100010011000101110001, 
24'b110100110010001011001111, 
24'b111110110101101110001110, 
24'b001011001111001011001111, 
24'b110111101111111100011011, 
24'b001011001111001011001111, 
24'b101000101001001010001111, 
24'b110100110001110100110001, 
24'b110110111111110001000000, 
24'b001011001111110100110001, 
24'b111100101010111110101101, 
24'b001011001111110100110001, 
24'b000010001000001100100101, 
24'b110100110001110100110001, 
24'b001111101110110100010011, 
24'b001011001111001011001111, 
24'b111110100100001001101000, 
24'b110100110001001011001111, 
24'b101101011100110001100010, 
24'b001011001111110100110001, 
24'b111011001100111111111010, 
24'b001011001111110100110001, 
24'b000001011010001111000111, 
24'b110100110001110100110001, 
24'b001110000010111110111000, 
24'b110100110001001011001111, 
24'b110100100011101111010011, 
24'b001011001111110100110001, 
24'b000010100010000101101100, 
24'b110100110001110100110001, 
24'b010001101011101101001110, 
24'b001011001111001011001111, 
24'b000001100100111001100011, 
24'b001011001111001011001111, 
24'b110010010011111110000110, 
24'b001011001111110100110001, 
24'b001001010000000010011111, 
24'b001011001111001011001111, 
24'b110001110011001110001001, 
24'b110100110001110100110001, 
24'b000000100001110011101110, 
24'b001011001111110100110001, 
24'b001111110111111111111010, 
24'b001011001111001011001111, 
24'b111111100010000110000001, 
24'b001011010000001011001111, 
24'b101111000000010100001000, 
24'b110100110010110100110001, 
24'b111101011011000100011101, 
24'b110100110001110100110001, 
24'b000100101011111100010101, 
24'b110100110001110100110001, 
24'b010011101001101100101001, 
24'b001011001111001011001111, 
24'b000101000000111010100111, 
24'b001011001111001011001111, 
24'b111110110100000000000100, 
24'b001011001111001011001111, 
24'b111000100001000101011101, 
24'b001011001111001011001111, 
24'b101001100000010011001001, 
24'b110100110001110100110000, 
24'b110111101000000010011100, 
24'b110100110001110100110000, 
24'b111100101110110010110011, 
24'b001011001111110100110001, 
24'b000000100100001001011001, 
24'b110100110001110100110001, 
24'b000101000100110001100010, 
24'b001011001111110100110001, 
24'b010001010100111111100010, 
24'b001011001111001011001111, 
24'b111000100000001101001110, 
24'b110100110001110100110001, 
24'b001101101010110011111000, 
24'b001011001111001011001111, 
24'b110101101111000001010010, 
24'b001011001111110100110001, 
24'b000111000001001100001010, 
24'b000000000000000000000000, 
24'b111101111100001011100100, 
24'b110100110001110100110001, 
24'b001000011111111111010010, 
24'b110100110001110100110001, 
24'b011000001100101111011100, 
24'b001011001111001011001111, 
24'b001010011000111110101010, 
24'b001011001111001011001111, 
24'b000101100101001100110010, 
24'b110100110001001011001111, 
24'b000010001110110011101011, 
24'b001011001111001011001111, 
24'b111111000000000001011010, 
24'b001011001111001011001111, 
24'b111010101001001111001011, 
24'b110100110001001011010000, 
24'b101101101101110110001101, 
24'b001011001111110100110001, 
24'b111111011001000100101000, 
24'b001011001111110100110001, 
24'b010001000100010100011101, 
24'b110100110001001011001111, 
24'b000100001001000101111001, 
24'b110100110010001011001111, 
24'b111111110001111111000101, 
24'b110100110001001011001111, 
24'b111100100010110001111100, 
24'b001011001111001011001111, 
24'b111001001010001010111011, 
24'b110100110001001011001111, 
24'b110100011001111100011000, 
24'b110100110001001011001111, 
24'b100110101100101100011101, 
24'b001011001111110100110001, 
24'b110110110110111010111111, 
24'b001011001111110100110000, 
24'b000101010110000001111110, 
24'b001011001111001011001111, 
24'b101100000001010000001010, 
24'b110100110001110100110001, 
24'b111000011110111111011000, 
24'b110100110010110100110001, 
24'b111110000011101110101101, 
24'b001011001111110100110001, 
24'b001001111111111101100010, 
24'b001011001111001011001111, 
24'b101111011000001011010010, 
24'b110100110001110100110001, 
24'b111010110001110001100110, 
24'b001011001111110100110001, 
24'b111110101001111101111110, 
24'b001011001111110100110001, 
24'b000001110101000011110011, 
24'b001011001111110100110001, 
24'b000101111101010000011110, 
24'b110100110001110100110001, 
24'b010010000000110111110110, 
24'b001011010000001011001111, 
24'b111001001001001101010000, 
24'b110100110001110100110000, 
24'b001110100001110110000010, 
24'b001011001111001011001111, 
24'b110111011100001011110100, 
24'b110100110001110100110001, 
24'b001101100110110100100101, 
24'b001011001111001011010000, 
24'b110111000111001001111011, 
24'b110100110001110100110001, 
24'b001110010111110001001101, 
24'b001011001111001011001111, 
24'b111111001101111101100110, 
24'b001011001111001011001111, 
24'b101111000101000010011111, 
24'b001011001111110100110001, 
24'b111101100111000111100101, 
24'b001011001111110100110001, 
24'b000100111001010101000110, 
24'b110100110001110100110001, 
24'b010011110000000100001010, 
24'b110100110010001011001111, 
24'b000100101110110011101101, 
24'b001011001111001011001111, 
24'b111101010000000011010101, 
24'b001011001111001011001110, 
24'b101110011111010011010010, 
24'b110100110000110100110001, 
24'b111110010101000100010111, 
24'b110100110001110100110001, 
24'b001100111111111100100111, 
24'b110100110001001011001111, 
24'b110100100001101101000011, 
24'b001011010000110100110001, 
24'b000011010000111010111110, 
24'b001011001111110100110001, 
24'b010011010000000000000000, 
24'b001011001111001011001111, 
24'b000100110100000011111101, 
24'b001011001111001011001111, 
24'b111110000010001000110011, 
24'b001011001111001011001111, 
24'b110000101110010110001011, 
24'b110100110000110100110001, 
24'b001000110110000101000010, 
24'b110100110001001011001111, 
24'b110010111110110100001010, 
24'b001011010000110100110001, 
24'b001001101101000010011010, 
24'b001011001111001011001111, 
24'b110011010101001001100100, 
24'b001011001111110100110001, 
24'b001001110001011000010110, 
24'b110100110001001011001111, 
24'b110011001001001000110100, 
24'b110100110001110100110001, 
24'b001001001101111010110110, 
24'b001011001111001011001111, 
24'b110001100100010100101011, 
24'b110100110000110100110001, 
24'b000000001111001000111100, 
24'b110100110001110100110001, 
24'b001111101001000101000100, 
24'b110100110001001011001111, 
24'b111111011100000010010000, 
24'b110100110000001011001111, 
24'b101111010000111111011011, 
24'b110100110001110100110001, 
24'b111110101011111011100110, 
24'b110100110001110100110001, 
24'b001101011011101111111101, 
24'b001011001111001011001111, 
24'b110110000001001001111000, 
24'b110100110001110100110001, 
24'b001101000000111100000011, 
24'b110100110001001011001111, 
24'b111101110001101100101101, 
24'b001011001111001011001111, 
24'b101101101101111011101101, 
24'b001011010000110100110001, 
24'b111100111010000011000101, 
24'b001011001111110100110001, 
24'b001011000000010001000011, 
24'b110100110001001011001111, 
24'b110001110101111001111101, 
24'b001011001111110100110001, 
24'b111111011010010001111011, 
24'b110100110001110100110001, 
24'b001100111011000100111101, 
24'b110100110001001011001111, 
24'b110011100000111111000100, 
24'b110100110001110100110001, 
24'b000001000100110010101111, 
24'b001011001110110100110001, 
24'b001110110001001100101100, 
24'b110100110001001011001111, 
24'b110110000010111111110111, 
24'b110100110001110100110001, 
24'b000111101111110110000110, 
24'b000000000000000000000000, 
24'b000011010000111011110100, 
24'b000000000000000000000000, 
24'b000010010100111101001110, 
24'b000000000000000000000000, 
24'b000001110111111101111010, 
24'b000000000000000000000000, 
24'b000001100110111110010110, 
24'b000000000000000000000000, 
24'b000001011010111110101000, 
24'b000000000000000000000000, 
24'b000001010000111110110110, 
24'b000000000000000000000000, 
24'b000001001000111111000000, 
24'b000000000000000000000000, 
24'b000001000011111111001000, 
24'b000000000001000000000000, 
24'b000000111110111111010000, 
24'b000000000000000000000000, 
24'b000000111001111111010101, 
24'b000000000000000000000000, 
24'b000000110110111111011010, 
24'b000000000000000000000000, 
24'b000000110011111111011101, 
24'b000000000000000000000000, 
24'b000000110000111111100001, 
24'b000000000000000000000000, 
24'b000000101110111111100100, 
24'b000000000000000000000000, 
24'b000000101100111111100111, 
24'b000000000000000000000000, 
24'b000000101010111111101001, 
24'b000000000000000000000000, 
24'b000000101000111111101100, 
24'b000000000000000000000000, 
24'b000000100111111111101101, 
24'b000000000000000000000000, 
24'b000000100101111111101111, 
24'b000000000000000000000000, 
24'b000000100100111111110001, 
24'b000000000000000000000000, 
24'b000000100011111111110010, 
24'b000000000000000000000000, 
24'b000000100010111111110011, 
24'b000000000000000000000000, 
24'b000000100000111111110100, 
24'b000000000000000000000000, 
24'b000000011111111111110110, 
24'b000000000000000000000000, 
24'b000000011110111111110111, 
24'b000000000000000000000000, 
24'b000000011110111111110111, 
24'b000000000000000000000000, 
24'b000000011101111111111000, 
24'b000000000000000000000000, 
24'b000000011100111111111001, 
24'b000000000000000000000000, 
24'b000000011100111111111010, 
24'b000000000000000000000000, 
24'b000000011011111111111010, 
24'b000000000000000000000000, 
24'b000000011010111111111011, 
24'b000000000000000000000000, 
24'b000000011010111111111011, 
24'b000000000000000000000000, 
24'b000000011001111111111100, 
24'b000000000000000000000000, 
24'b000000011001111111111101, 
24'b000000000000000000000000, 
24'b000000011000111111111101, 
24'b000000000000000000000000, 
24'b000000011000111111111101, 
24'b000000000000000000000000, 
24'b000000010111111111111110, 
24'b000000000000000000000000, 
24'b000000010111111111111110, 
24'b000000000000000000000000, 
24'b000000010110111111111111, 
24'b000000000000000000000000, 
24'b000000010110111111111111, 
24'b000000000000000000000000, 
24'b000000010101111111111111, 
24'b000000000000000000000000, 
24'b000000010101111111111111, 
24'b000000000000000000000000, 
24'b000000010101111111111111, 
24'b000000000000000000000000, 
24'b000000010100000000000000, 
24'b000000000000000000000000, 
24'b000000010100000000000000, 
24'b000000000000000000000000, 
24'b000000010100000000000000, 
24'b000000000000000000000000, 
24'b000000010011000000000001, 
24'b000000000000000000000000, 
24'b000000010011000000000000, 
24'b000000000000000000000000, 
24'b000000010011000000000001, 
24'b000000000000000000000000, 
24'b000000010011000000000001, 
24'b000000000000000000000000, 
24'b000000010011000000000001, 
24'b000000000000000000000000, 
24'b000000010011000000000010, 
24'b000000000000000000000001, 
24'b000000010001000000000001, 
24'b000000000000000000000000, 
24'b000000010010000000000010, 
24'b000000000000000000000000, 
24'b000000010001000000000010, 
24'b000000000000000000000000, 
24'b000000010001000000000010, 
24'b000000000000000000000000, 
24'b000000010001000000000010, 
24'b000000000000000000000000, 
24'b000000010001000000000010, 
24'b000000000000000000000000, 
24'b000000010001000000000011, 
24'b000000000000000000000000, 
24'b000000010001000000000010, 
24'b000000000000000000000001, 
24'b000000010000000000000010, 
24'b000000000000000000000000, 
24'b000000010000000000000010, 
24'b000000000000000000000000, 
24'b000000001111000000000011, 
24'b000000000000000000000000, 
24'b000000010000000000000010, 
24'b000000000000000000000000, 
24'b000000010000000000000011, 
24'b000000000000000000000000, 
24'b000000001111000000000011, 
24'b000000000000000000000000, 
24'b000000001111000000000011, 
24'b000000000000111111111111, 
24'b000000001111000000000011, 
24'b000000000000000000000000, 
24'b000000001111000000000011, 
24'b000000000000000000000000, 
24'b000000001111000000000011, 
24'b000000000000000000000000, 
24'b000000001111000000000011, 
24'b000000000000000000000000, 
24'b000000001110000000000011, 
24'b000000000000000000000000, 
24'b000000001111000000000011, 
24'b000000000000000000000000, 
24'b000000001110000000000011, 
24'b000000000000000000000000, 
24'b000000001110000000000011, 
24'b000000000000000000000000, 
24'b000000001110000000000011, 
24'b000000000000000000000000, 
24'b000000001110000000000011, 
24'b000000000000000000000000, 
24'b000000001110000000000011, 
24'b000000000000000000000000, 
24'b000000001110000000000011, 
24'b000000000000000000000001, 
24'b000000001101000000000011, 
24'b000000000000000000000000, 
24'b000000001101000000000011, 
24'b000000000000000000000000, 
24'b000000001101000000000011, 
24'b000000000000000000000000, 
24'b000000001101000000000100, 
24'b000000000000000000000000, 
24'b000000001101000000000011, 
24'b000000000000000000000000, 
24'b000000001101000000000100, 
24'b000000000000000000000000, 
24'b000000001101000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000000000000000000, 
24'b000000001101000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000011, 
24'b000000000001000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001100000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000001, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001011000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b111111111111000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000001, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000001000000000000, 
24'b000000001010000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000111111111111, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000100, 
24'b000000000000000000000000, 
24'b000000001010000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000111111111111, 
24'b000000001010000000000011, 
24'b000000000000000000000001, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000010, 
24'b000000000001000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000010, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000011, 
24'b000000000000000000000001, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001001000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000111111111111, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000011, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000001, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000001, 
24'b000000000000000000000001, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000001000000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000001000000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000010, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000111111111111, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000001000000000000001, 
24'b000000000000000000000000, 
24'b000000001000000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000001, 
24'b000000000000111111111111, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000111111111111, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000001000000000000, 
24'b000000000111000000000001, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000111111111111, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000001, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000001, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111000000000000, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000001000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000001000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110000000000000, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000000, 
24'b000000000111111111111111, 
24'b000000000000000000000001, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b000000000110111111111111, 
24'b000000000000000000000000, 
24'b0_00000000111111111111110, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000100, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000001000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000010000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000011000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000110, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000110, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000110, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000110, 
24'b000000000000000000000000, 
24'b000000000100000000000110, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000000000000000001, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000100000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000111111111111, 
24'b000000000110000000000110, 
24'b000000000000000000000001, 
24'b000000000101000000000101, 
24'b000000000000000000000000, 
24'b000000000101000000000101, 
24'b000000000001000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000101000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000110000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000000111000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001000000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001001000000000111, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000111, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000111, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000111, 
24'b000000000000000000000000, 
24'b000000001010000000000111, 
24'b000000000000000000000000, 
24'b000000001010000000000110, 
24'b000000000000000000000000, 
24'b000000001010000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001010000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001011000000000111, 
24'b000000000000000000000000, 
24'b000000001100000000000111, 
24'b000000000000000000000000, 
24'b000000001100000000000111, 
24'b000000000000000000000000, 
24'b000000001100000000000111, 
24'b000000000000000000000000, 
24'b000000001100000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001100000000000111, 
24'b000000000000000000000000, 
24'b000000001100000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001101000000000111, 
24'b000000000000000000000000, 
24'b000000001110000000000111, 
24'b000000000000000000000000, 
24'b000000001110000000000111, 
24'b000000000000000000000000, 
24'b000000001110000000000111, 
24'b000000000000000000000000, 
24'b000000001110000000000111, 
24'b000000000000000000000000, 
24'b000000001111000000000111, 
24'b000000000000000000000000, 
24'b000000001110000000000111, 
24'b000000000000000000000000, 
24'b000000001110000000000111, 
24'b000000000000000000000000, 
24'b000000001111000000001000, 
24'b000000000000000000000000, 
24'b000000001111000000001000, 
24'b000000000000000000000000, 
24'b000000001111000000000111, 
24'b000000000000000000000000, 
24'b000000001111000000000111, 
24'b000000000000000000000000, 
24'b000000010000000000000111, 
24'b000000000000000000000000, 
24'b000000010000000000000111, 
24'b000000000000000000000000, 
24'b000000010000000000001000, 
24'b000000000000000000000000, 
24'b000000010000000000001000, 
24'b000000000000000000000000, 
24'b000000010000000000001000, 
24'b000000000000000000000000, 
24'b000000010000000000001000, 
24'b000000000000000000000000, 
24'b000000010001000000000111, 
24'b000000000000000000000000, 
24'b000000010001000000001000, 
24'b000000000000000000000000, 
24'b000000010010000000001000, 
24'b000000000000000000000000, 
24'b000000010010000000001000, 
24'b000000000000000000000000, 
24'b000000010010000000001000, 
24'b000000000000000000000000, 
24'b000000010010000000001000, 
24'b000000000000000000000000, 
24'b000000010010000000001000, 
24'b000000000000000000000000, 
24'b000000010011000000001000, 
24'b000000000000000000000000, 
24'b000000010011000000001000, 
24'b000000000000000000000000, 
24'b000000010011000000001000, 
24'b000000000000000000000000, 
24'b000000010011000000001000, 
24'b000000000000000000000000, 
24'b000000010100000000001000, 
24'b000000000000000000000000, 
24'b000000010100000000001000, 
24'b000000000000000000000000, 
24'b000000010100000000001001, 
24'b000000000000000000000000, 
24'b000000010101000000001001, 
24'b000000000000000000000000, 
24'b000000010101000000001000, 
24'b000000000000000000000000, 
24'b000000010101000000001000, 
24'b000000000000000000000000, 
24'b000000010101000000001001, 
24'b000000000000000000000000, 
24'b000000010110000000001001, 
24'b000000000000000000000000, 
24'b000000010111000000001000, 
24'b000000000000000000000000, 
24'b000000010111000000001001, 
24'b000000000000000000000000, 
24'b000000010111000000001001, 
24'b000000000000000000000000, 
24'b000000011000000000001001, 
24'b000000000000000000000000, 
24'b000000011000000000001001, 
24'b000000000000000000000000, 
24'b000000011000000000001001, 
24'b000000000000000000000000, 
24'b000000011001000000001001, 
24'b000000000000000000000000, 
24'b000000011001000000001001, 
24'b000000000000000000000000, 
24'b000000011010000000001001, 
24'b000000000000000000000000, 
24'b000000011011000000001001, 
24'b000000000000000000000000, 
24'b000000011011000000001001, 
24'b000000000000000000000000, 
24'b000000011011000000001010, 
24'b000000000000000000000000, 
24'b000000011100000000001001, 
24'b000000000000000000000000, 
24'b000000011101000000001010, 
24'b000000000000000000000000, 
24'b000000011101000000001001, 
24'b000000000000000000000000, 
24'b000000011110000000001010, 
24'b000000000000000000000000, 
24'b000000011110000000001010, 
24'b000000000000000000000000, 
24'b000000011111000000001010, 
24'b000000000000000000000000, 
24'b000000100000000000001010, 
24'b000000000000000000000000, 
24'b000000100001000000001010, 
24'b000000000000000000000000, 
24'b000000100010000000001010, 
24'b000000000000000000000000, 
24'b000000100010000000001010, 
24'b000000000000000000000000, 
24'b000000100011000000001010, 
24'b000000000000000000000000, 
24'b000000100100000000001010, 
24'b000000000000000000000000, 
24'b000000100101000000001011, 
24'b000000000000000000000000, 
24'b000000100101000000001011, 
24'b000000000000000000000000, 
24'b000000100111000000001010, 
24'b000000000000000000000000, 
24'b000000101000000000001011, 
24'b000000000000000000000000, 
24'b000000101001000000001011, 
24'b000000000000000000000000, 
24'b000000101010000000001011, 
24'b000000000000000000000000, 
24'b000000101011000000001011, 
24'b000000000000000000000000, 
24'b000000101101000000001011, 
24'b000000000000000000000000, 
24'b000000101110000000001011, 
24'b000000000000000000000000, 
24'b000000110000000000001011, 
24'b000000000000000000000000, 
24'b000000110010000000001100, 
24'b000000000000000000000000, 
24'b000000110011000000001100, 
24'b000000000000000000000000, 
24'b000000110101000000001011, 
24'b000000000000000000000000, 
24'b000000110111000000001011, 
24'b000000000000000000000000, 
24'b000000111001000000001100, 
24'b000000000000000000000000, 
24'b000000111011000000001011, 
24'b000000000000000000000000, 
24'b000000111110000000001011, 
24'b000000000000000000000000, 
24'b000001000001000000001011, 
24'b000000000000000000000000, 
24'b000001000100000000001011, 
24'b000000000000000000000000, 
24'b000001000111000000001011, 
24'b000000000000000000000000, 
24'b000001001010000000001011, 
24'b000000000000000000000000, 
24'b000001001110000000001010, 
24'b000000000000000000000000, 
24'b000001010010000000001010, 
24'b000000000000000000000000, 
24'b000001010111000000001000, 
24'b000000000000000000000000, 
24'b000001011100000000001000, 
24'b000000000000000000000000, 
24'b000001100010000000000111, 
24'b000000000000000000000000, 
24'b000001101001000000000100, 
24'b000000000000000000000000, 
24'b000001110001000000000010, 
24'b000000000000000000000000, 
24'b000001111001111111111110, 
24'b000000000000000000000000, 
24'b000010000011111111111001, 
24'b000000000000000000000000, 
24'b000010001110111111110001, 
24'b000000000000000000000000, 
24'b000010011100111111100101, 
24'b000000000000000000000000, 
24'b000010101011111111010001, 
24'b000000000000000000000000, 
24'b000010111001111110101010, 
24'b000000000000000000000000, 
24'b000010110111111101001111, 
24'b000000000000000000000000, 
24'b111111000111110110100110, 
24'b001101111100110010000100, 
24'b011000101101000011011010, 
24'b001101111100001101111100, 
24'b001000011000010100011110, 
24'b110010000100001101111100, 
24'b000001010010110110110010, 
24'b001101111100001101111100, 
24'b110010011110010010000110, 
24'b110010000100110010000100, 
24'b010011100110110110001001, 
24'b001101111100001101111100, 
24'b000101100110010010010010, 
24'b110010000100001101111100, 
24'b000000111111110111001100, 
24'b001101111100001101111100, 
24'b111101010010010101000010, 
24'b110010000100001101111100, 
24'b111000100101000011110101, 
24'b110010000011001101111100, 
24'b101010010111110011001001, 
24'b001101111100110010000100, 
24'b001010111111010011010000, 
24'b110010000100001101111100, 
24'b111010110010000100010001, 
24'b110010000100001101111100, 
24'b101010001011111110010100, 
24'b110010000100110010000100, 
24'b001001011010110111110111, 
24'b110010000100001101111100, 
24'b110111101001100110101010, 
24'b001101111100001101111100, 
24'b100011111110111010001001, 
24'b001101111100110010000100, 
24'b110101101101000100001111, 
24'b001101111100110010000100, 
24'b111100111011010111101101, 
24'b110010000100110010000100, 
24'b000100000010000110011011, 
24'b110010000100110010000100, 
24'b010101010101111111110101, 
24'b110010000100001101111100, 
24'b000000101100111001101011, 
24'b110010000100001101111100, 
24'b101100011111101010010111, 
24'b001101111100110010000100, 
24'b111111101111001001111100, 
24'b110010000100110010000100, 
24'b010010010100111000010010, 
24'b110010000100001101111100, 
24'b110101101100100100110011, 
24'b001101111100110010000100, 
24'b010010100111110111001010, 
24'b001101111100001101111100, 
24'b111101001100000011010011, 
24'b000000000000000000000000, 
24'b001001010000110110010111, 
24'b001101111100001101111100, 
24'b111110100100000001111011, 
24'b001101111100001101111100, 
24'b110111001101010010011101, 
24'b110010000100001101111100, 
24'b100101011110110100011001, 
24'b001101111100110010000100, 
24'b111000011111001111011001, 
24'b110010000100110010000100, 
24'b000001111101110011000100, 
24'b001101111100110010000100, 
24'b010100011010001110101110, 
24'b110010000100001101111100, 
24'b000000110001110010110001, 
24'b001101111101001101111100, 
24'b101110011000001110110001, 
24'b110010000100110010000100, 
24'b001011101110110011010011, 
24'b001101111100001101111100, 
24'b110000100001010000100111, 
24'b110010000100110010000100, 
24'b001100111100111110100001, 
24'b110010000100001101111100, 
24'b110001111010101100010010, 
24'b001101111100110010000100, 
24'b001111110011001001000010, 
24'b110010000100001101111100, 
24'b111111001000101011111000, 
24'b001101111100001101111100, 
24'b110110010111111101100110, 
24'b001101111100001101111100, 
24'b100011101100001110111000, 
24'b110010000100110010000100, 
24'b110101100010101111101101, 
24'b001101111100110010000100, 
24'b111100101001000000110110, 
24'b001101111100110010000011, 
24'b000011100000010010001111, 
24'b110010000100110010000100, 
24'b010100011110110100010111, 
24'b001101111100001101111100, 
24'b111111010110001111000101, 
24'b110010000100001101111100, 
24'b101010010100110001100011, 
24'b001101111100110010000100, 
24'b111011101100000011111000, 
24'b001101111100110010000011, 
24'b000011111111010111011110, 
24'b110010000100110010000101, 
24'b010101000000000100110000, 
24'b110010000100001101111100, 
24'b111011111001110111010011, 
24'b000000000000000000000000, 
24'b111111111110111101101000, 
24'b000000000000000000000000, 
24'b000000010011111110111000, 
24'b000000000000000000000000, 
24'b000000010010111111010111, 
24'b000000000000000000000000, 
24'b000000001110111111100110, 
24'b000000000000000000000000, 
24'b000000001010111111110000, 
24'b000000000000000000000000, 
24'b000000000111111111110101, 
24'b000000000000000000000000, 
24'b000000000100111111111000, 
24'b000000000000000000000000, 
24'b000000000001111111111011, 
24'b000000000000000000000000, 
24'b111111111111111111111101, 
24'b000000000000000000000000, 
24'b111111111101111111111110, 
24'b000000000000000000000000, 
24'b111111111100111111111111, 
24'b000000000000000000000000, 
24'b111111111010111111111111, 
24'b000000000000000000000000, 
24'b111111111001000000000000, 
24'b000000000000000000000000, 
24'b111111111000000000000000, 
24'b000000000000000000000000, 
24'b111111111000000000000001, 
24'b000000000000000000000000, 
24'b111111110111000000000001, 
24'b000000000000111111111111, 
24'b111111110111000000000001, 
24'b000000000000000000000000, 
24'b111111110110000000000001, 
24'b000000000000000000000000, 
24'b111111110110000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110011000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110011000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110011000000000010, 
24'b000000000000000000000000, 
24'b111111110011000000000010, 
24'b000000000000000000000000, 
24'b111111110011000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110011000000000010, 
24'b000000000000000000000000, 
24'b111111110011000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000010, 
24'b000000000000000000000000, 
24'b111111110100000000000011, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110101000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000010, 
24'b000000000000000000000000, 
24'b111111110101000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000010, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000010, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000010, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110110000000000010, 
24'b000000000000000000000000, 
24'b111111110110000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111110111000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111000000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111001000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111010000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111010000000000100, 
24'b000000000000111111111111, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000111111111111, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111011000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b111111111111000000000000, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000011, 
24'b000000000000000000000000, 
24'b111111111101000000000011, 
24'b000000000000000000000000, 
24'b111111111100000000000011, 
24'b000000000001000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111100000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111101000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111110000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000100, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b000000000000000000000101, 
24'b000000000000000000000000, 
24'b111111111111000000000101, 
24'b000000000000000000000000, 
24'b0_00000000000000000000101, 
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b111111111111000000000000,
24'b000000000011000000000111,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001010000000001011,
24'b000000000000000000000000,
24'b000000001010000000001011,
24'b000000000000000000000000,
24'b000000001010000000001011,
24'b000000000000000000000000,
24'b000000001010000000001100,
24'b000000000000000000000000,
24'b000000001010000000001100,
24'b000000000000000000000000,
24'b000000001010000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001101,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001101,
24'b000000000000000000000000,
24'b000000001100000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000010000000000001110,
24'b000000000000000000000000,
24'b000000010000000000001110,
24'b000000000000000000000000,
24'b000000010000000000001110,
24'b000000000000000000000000,
24'b000000010001000000001110,
24'b000000000000000000000000,
24'b000000010001000000001110,
24'b000000000000000000000000,
24'b000000010001000000001111,
24'b000000000000000000000000,
24'b000000010001000000001111,
24'b000000000000000000000000,
24'b000000010010000000001111,
24'b000000000000000000000000,
24'b000000010010000000001111,
24'b000000000000000000000000,
24'b000000010010000000001111,
24'b000000000000000000000000,
24'b000000010011000000001111,
24'b000000000000000000000000,
24'b000000010011000000001111,
24'b000000000000000000000000,
24'b000000010011000000001111,
24'b000000000000000000000000,
24'b000000010100000000010000,
24'b000000000000000000000000,
24'b000000010100000000010000,
24'b000000000000000000000000,
24'b000000010100000000010000,
24'b000000000000000000000000,
24'b000000010101000000010000,
24'b000000000000000000000000,
24'b000000010101000000010000,
24'b000000000000000000000000,
24'b000000010110000000010000,
24'b000000000000000000000000,
24'b000000010110000000010000,
24'b000000000000000000000000,
24'b000000010110000000010000,
24'b000000000000000000000000,
24'b000000010111000000010001,
24'b000000000000000000000000,
24'b000000010111000000010001,
24'b000000000000000000000000,
24'b000000010111000000010001,
24'b000000000000000000000000,
24'b000000011000000000010001,
24'b000000000000000000000000,
24'b000000011000000000010001,
24'b000000000000000000000000,
24'b000000011001000000010001,
24'b000000000000000000000000,
24'b000000011001000000010010,
24'b000000000000000000000000,
24'b000000011010000000010010,
24'b000000000000000000000000,
24'b000000011011000000010010,
24'b000000000000000000000000,
24'b000000011011000000010010,
24'b000000000000000000000000,
24'b000000011100000000010010,
24'b000000000000000000000000,
24'b000000011100000000010010,
24'b000000000000000000000000,
24'b000000011101000000010011,
24'b000000000000000000000000,
24'b000000011101000000010011,
24'b000000000000000000000000,
24'b000000011110000000010011,
24'b000000000000000000000000,
24'b000000011111000000010011,
24'b000000000000000000000000,
24'b000000100000000000010100,
24'b000000000000000000000000,
24'b000000100000000000010100,
24'b000000000000000000000000,
24'b000000100001000000010100,
24'b000000000000000000000000,
24'b000000100010000000010100,
24'b000000000000000000000000,
24'b000000100011000000010100,
24'b000000000000000000000000,
24'b000000100100000000010101,
24'b000000000000000000000000,
24'b000000100101000000010101,
24'b000000000000000000000000,
24'b000000100110000000010101,
24'b000000000000000000000000,
24'b000000100111000000010101,
24'b000000000000000000000000,
24'b000000101000000000010101,
24'b000000000000000000000000,
24'b000000101001000000010110,
24'b000000000000000000000000,
24'b000000101011000000010110,
24'b000000000000000000000000,
24'b000000101100000000010110,
24'b000000000000000000000000,
24'b000000101101000000010111,
24'b000000000000000000000000,
24'b000000101111000000010111,
24'b000000000000000000000000,
24'b000000110001000000010111,
24'b000000000000000000000000,
24'b000000110010000000011000,
24'b000000000000000000000000,
24'b000000110100000000011000,
24'b000000000000000000000000,
24'b000000110110000000011000,
24'b000000000000000000000000,
24'b000000111000000000011000,
24'b000000000000000000000000,
24'b000000111010000000011000,
24'b000000000000000000000000,
24'b000000111101000000011001,
24'b000000000000000000000000,
24'b000001000000000000011001,
24'b000000000000000000000000,
24'b000001000010000000011001,
24'b000000000000000000000000,
24'b000001000110000000011001,
24'b000000000000000000000000,
24'b000001001001000000011001,
24'b000000000000000000000000,
24'b000001001100000000011001,
24'b000000000000000000000000,
24'b000001010001000000011001,
24'b000000000000000000000000,
24'b000001010101000000011001,
24'b000000000000000000000000,
24'b000001011010000000011000,
24'b000000000000000000000000,
24'b000001100000000000010111,
24'b000000000000000000000000,
24'b000001100110000000010110,
24'b000000000000000000000000,
24'b000001101101000000010100,
24'b000000000000000000000000,
24'b000001110110000000010010,
24'b000000000000000000000000,
24'b000001111111000000001110,
24'b000000000000000000000000,
24'b000010001010000000001001,
24'b000000000000000000000000,
24'b000010010111000000000000,
24'b000000000000000000000000,
24'b000010100101111111110100,
24'b000000000000000000000000,
24'b000010110110111111011101,
24'b000000000000000000000000,
24'b000011000101111110110011,
24'b000000000000000000000000,
24'b000011000010111101001111,
24'b000000000000000000000000,
24'b111110110111110101110110,
24'b001111011111110000100001,
24'b011011010010000100000110,
24'b001111011111001111011111,
24'b001001001001010111000100,
24'b110000100001001111011111,
24'b000001001111110110000101,
24'b001111011111001111011111,
24'b110000110010010100011011,
24'b110000100001110000100001,
24'b010101100101110101011001,
24'b001111011111001111011111,
24'b000110000000010100101100,
24'b110000100001001111011110,
24'b000000110111110110100101,
24'b001111011111001111011111,
24'b111100101110010111110000,
24'b110000100001001111011111,
24'b110111011101000100101010,
24'b110000100001001111011111,
24'b100111100110110010001000,
24'b001111011111110000100001,
24'b001011101111010101110010,
24'b110000100001001111011111,
24'b111001011110000101000101,
24'b110000100001001111011111,
24'b100110001110111110000101,
24'b110000100001110000100001,
24'b000011010100110010101010,
24'b000000000000000000000000,
24'b000101101100111111111010,
24'b110000100001001111011111,
24'b110110001000100110100110,
24'b001111011111001111011111,
24'b100000100110111011001110,
24'b001111011111110000100001,
24'b110100010010000110000011,
24'b001111011111110000100001,
24'b111100001111011011100010,
24'b110000100001110000100001,
24'b000100000010001000010010,
24'b110000100001110000100001,
24'b010111001000000000111110,
24'b110000100001001111011111,
24'b000000000101111010001011,
24'b110000100010001111011111,
24'b101001011101101001010100,
24'b001111011111110000100001,
24'b111110101000001100100011,
24'b110000100001110000100001,
24'b010010111100111001001100,
24'b110000100010001111011111,
24'b110010101001100011111110,
24'b001111011111110000100001,
24'b010001111100111001000110,
24'b001111011111001111011111,
24'b111000010010001000010001,
24'b000000000000000000000000,
24'b111101101110000001011001,
24'b000000000000000000000000,
24'b111110100011000000001001,
24'b000000000000000000000000,
24'b111110110110111111101101,
24'b000000000000000000000000,
24'b111110111111111111100010,
24'b000000000000000000000000,
24'b111111000101111111011100,
24'b000000000000000000000000,
24'b111111001000111111011010,
24'b000000000000000000000000,
24'b111111001011111111011010,
24'b000000000000000000000000,
24'b111111001101111111011010,
24'b000000000000000000000000,
24'b111111001111111111011011,
24'b000000000000000000000000,
24'b111111010000111111011100,
24'b000000000000000000000000,
24'b111111010010111111011101,
24'b000000000000000000000000,
24'b111111010011111111011110,
24'b000000000000000000000000,
24'b111111010100111111011111,
24'b000000000000000000000000,
24'b111111010101111111100000,
24'b000000000000000000000000,
24'b111111010110111111100001,
24'b000000000000000000000000,
24'b111111010111111111100010,
24'b000000000000000000000000,
24'b111111011000111111100100,
24'b000000000000000000000000,
24'b111111011001111111100101,
24'b000000000000000000000000,
24'b111111011010111111100110,
24'b000000000000000000000000,
24'b111111011011111111100110,
24'b000000000000000000000000,
24'b111111011011111111100111,
24'b000000000000000000000000,
24'b111111011100111111101000,
24'b000000000000000000000000,
24'b111111011101111111101001,
24'b000000000000000000000000,
24'b111111011110111111101010,
24'b000000000000000000000000,
24'b111111011110111111101010,
24'b000000000000000000000000,
24'b111111011111111111101011,
24'b000000000000000000000000,
24'b111111011111111111101100,
24'b000000000000000000000000,
24'b111111100000111111101100,
24'b000000000000000000000000,
24'b111111100000111111101101,
24'b000000000000000000000000,
24'b111111100001111111101110,
24'b000000000000000000000000,
24'b111111100001111111101110,
24'b000000000000000000000000,
24'b111111100010111111101111,
24'b000000000000000000000000,
24'b111111100010111111101111,
24'b000000000000000000000000,
24'b111111100011111111101111,
24'b000000000000000000000000,
24'b111111100011111111110000,
24'b000000000000000000000000,
24'b111111100100111111110000,
24'b000000000000000000000000,
24'b111111100100111111110001,
24'b000000000000000000000000,
24'b111111100100111111110001,
24'b000000000000000000000000,
24'b111111100101111111110010,
24'b000000000000000000000000,
24'b111111100101111111110010,
24'b000000000000000000000000,
24'b111111100101111111110011,
24'b000000000000000000000000,
24'b111111100110111111110011,
24'b000000000000000000000000,
24'b111111100110111111110011,
24'b000000000000000000000000,
24'b111111100111111111110011,
24'b000000000000000000000000,
24'b111111100111111111110100,
24'b000000000000000000000000,
24'b111111100111111111110100,
24'b000000000000000000000000,
24'b111111101000111111110100,
24'b000000000000000000000000,
24'b111111101000111111110101,
24'b000000000000000000000000,
24'b111111101000111111110101,
24'b000000000000000000000000,
24'b111111101000111111110101,
24'b000000000000000000000000,
24'b111111101001111111110101,
24'b000000000000000000000000,
24'b111111101001111111110110,
24'b000000000000000000000000,
24'b111111101010111111110110,
24'b000000000000000000000000,
24'b111111101001111111110110,
24'b000000000000000000000000,
24'b111111101010111111110110,
24'b000000000000000000000000,
24'b111111101010111111110111,
24'b000000000000000000000000,
24'b111111101010111111110111,
24'b000000000000000000000000,
24'b111111101010111111110111,
24'b000000000000000000000000,
24'b111111101011111111110111,
24'b000000000000000000000000,
24'b111111101011111111110111,
24'b000000000000000000000000,
24'b111111101011111111111000,
24'b000000000000000000000000,
24'b111111101011111111111000,
24'b000000000000000000000000,
24'b111111101100111111111000,
24'b000000000000000000000000,
24'b111111101100111111111000,
24'b000000000000000000000000,
24'b111111101100111111111000,
24'b000000000000000000000000,
24'b111111101100111111111001,
24'b000000000000000000000000,
24'b111111101100111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111010,
24'b000000000000000000000000,
24'b111111101101111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111110000111111111011,
24'b000000000000000000000000,
24'b111111110000111111111011,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111101,
24'b000000000000000000000000,
24'b111111110011111111111101,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110111000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101};