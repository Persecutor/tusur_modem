logic [23:0]	rom_freq_pr [0:1023] = {
24'b111000011001001000110101,
24'b000111101001111010100000,
24'b111101000100111000100000,
24'b000101110001001011100110,
24'b111101100010110011001011,
24'b111000010100001111100101,
24'b001000010001110111000111,
24'b111011100011111110111011,
24'b000100010001000010010011,
24'b000001100000111111100010,
24'b111000100111111110110111,
24'b000001011001000011011110,
24'b000001111100000010011011,
24'b000101111101110011001011,
24'b111100001100001010101000,
24'b110011110111111110010100,
24'b010000101000000010100100,
24'b111011100000111011001111,
24'b111101000000111101110101,
24'b111100110101000011000101,
24'b001100100100001100110011,
24'b110001001111100101110101,
24'b001001100111010000011110,
24'b111100101100000011101001,
24'b111111101101111000111100,
24'b000001111100111100011011,
24'b111111100110000100011000,
24'b111010000001000011100011,
24'b001100110000111111101000,
24'b110011011011110101101000,
24'b000100100000001010100001,
24'b000011100111111111111001,
24'b111010101111111001110000,
24'b000011010101111111001101,
24'b111111011000001101000000,
24'b111100111110110111000111,
24'b111111110101110101101111,
24'b001010001101001101101000,
24'b111001110110000010011011,
24'b110101010101111010000000,
24'b000111001011111011110101,
24'b001100000010000010001011,
24'b110110011001000011100101,
24'b111101001110000110011011,
24'b111011111000110001110110,
24'b000101100000000100000101,
24'b001111001101000101010000,
24'b101011100111111100000100,
24'b000001011011000011110100,
24'b000110011101111011100010,
24'b111111110011111101110110,
24'b111100001011001001101011,
24'b001010101011110110011111,
24'b110001100000000100011001,
24'b000011000010111111011111,
24'b000110000101000000111100,
24'b111110000111111101000001,
24'b000011010011000001110000,
24'b110110011111111111001001,
24'b000000100011000101101001,
24'b001101110110110111001001,
24'b110111100001000011100111,
24'b110011101110000010101111,
24'b010101000110111011111111,
24'b110111011000000011011111,
24'b111101001001111101010010,
24'b111110101100000011001001,
24'b000100101010110111010010,
24'b111111000010001101100111,
24'b000011111010110111100010,
24'b111011100100111111101110,
24'b111010010100000000101000,
24'b000010110011000101101010,
24'b001011000101110110000010,
24'b111000101100001000010010,
24'b000001000100111100101011,
24'b110110110001000010100010,
24'b000001101001111100000011,
24'b010000100101111101001111,
24'b111001011000001001001010,
24'b111001001001000000011110,
24'b111000001001110111001001,
24'b001111010111111010111101,
24'b111100110000010001100000,
24'b000011100100111010011100,
24'b111001111000111001101110,
24'b111001110010111110001001,
24'b001001101000001011001011,
24'b111100110001110110011010,
24'b000011100001000111001001,
24'b000100001000111011000000,
24'b110001010110111110001010,
24'b000100100100000110110100,
24'b000010101001111111111111,
24'b001001101100110001010001,
24'b110110010001010001000110,
24'b111110011100000001011011,
24'b111100000110110010111101,
24'b001010001101111111010011,
24'b111011100100001010001001,
24'b000101111101000000101101,
24'b110111101110111101110110,
24'b111111000111110111001011,
24'b000011010000000011101001,
24'b000000111000000111001101,
24'b000011110100111110110100,
24'b111011110010111011011000,
24'b111100100111000001111111,
24'b000001110101111010001010,
24'b000001011011000110010001,
24'b000010111110000011010010,
24'b111101111001000001110000,
24'b111111110011101110101101,
24'b111010101011001110001100,
24'b000101010101111100111101,
24'b000000100001000011010110,
24'b000000100011111111111100,
24'b111111100010110110001011,
24'b111011100000001000111011,
24'b000100111101111101100000,
24'b111000110001000001010100,
24'b001011010111111111011000,
24'b111100010010000010010010,
24'b111100101000111001111110,
24'b111011011000000001010101,
24'b001011100101000101001111,
24'b110101011000111100111011,
24'b001010011000000010010010,
24'b111000111101111010000100,
24'b000100001011000111010111,
24'b111000110000110011111101,
24'b000001111101001101111011,
24'b000100000101111110000111,
24'b001010010011111100101010,
24'b101100011110111010110001,
24'b000101000000111101101000,
24'b000000001101010000100000,
24'b000011100000111100001011,
24'b001101110010111000000101,
24'b100111000101111011000000,
24'b000110111101000010011000,
24'b000001111001010010100001,
24'b000101011011110011010011,
24'b000000110100111100110111,
24'b111001010011111010101111,
24'b000000100110000111101101,
24'b111000111011001000100111,
24'b001110001110110111010110,
24'b000001101100000000001100,
24'b110110000101110110111111,
24'b111100011010001001010101,
24'b000000100001001100111010,
24'b010010011011101000111000,
24'b110011100100001001111011,
24'b110110010101000100000000,
24'b001000100111110111101100,
24'b001000101100000011011101,
24'b110101111011000110000010,
24'b000010000000111000001110,
24'b110101101100000010111111,
24'b010101111010111101000110,
24'b110101100010000100101100,
24'b111010010100111011110110,
24'b000011001110000100111100,
24'b111111110111111010111101,
24'b000100100100000101011010,
24'b111110100000110111000000,
24'b000010011101000101011110,
24'b110100001001000011011011,
24'b000000010110000011010010,
24'b010011111110101111000101,
24'b111000101101001010111011,
24'b101111010001000001100110,
24'b001101000001000010010101,
24'b111111101010110111111001,
24'b111101111011000010011010,
24'b000110000000000001101000,
24'b110100111101000000011010,
24'b001011101000000000011010,
24'b111000100010111011101011,
24'b111000101011000111011001,
24'b010000111100111001100001,
24'b111100110001000000000110,
24'b111010001011000100011101,
24'b111011001011111101111110,
24'b000100101101000001011111,
24'b000010100011111000100101,
24'b000100001011001001101011,
24'b000001100101111110100010,
24'b101100110000111001010011,
24'b000100110010000000001111,
24'b010100100000001010100101,
24'b110100100000111111110001,
24'b111110001101101101100111,
24'b111010101111001010011010,
24'b000011101011000101011001,
24'b000110001010000101001011,
24'b111001100010110101010111,
24'b001011100111110010100101,
24'b101110001111010100110101,
24'b000101111111111111001101,
24'b000111000010000011101111,
24'b110110011110101010111111,
24'b001100111001000111111011,
24'b110110100101001000110101,
24'b111110110110000100000010,
24'b000000000100110011110011,
24'b000010100100111101011010,
24'b000000111101001010101101,
24'b001011110111111001011000,
24'b100110000010000100110010,
24'b001001010111111110111001,
24'b001000111101111011110100,
24'b111100001110000100011001,
24'b000100010010111011001101,
24'b110100000011000011100101,
24'b000010101000000100100000,
24'b000101010001111000101111,
24'b000001100001000010101001,
24'b000001011110111010011011,
24'b110100001110001011100000,
24'b000111100111110110101011,
24'b000000000111000110110111,
24'b000001011111111011111011,
24'b111101100011111011011001,
24'b111110001100000100110101,
24'b000111001011000100100001,
24'b111000001001111110100101,
24'b000000011010111001010110,
24'b000000011000111101111011,
24'b001101111011001011001100,
24'b101110100000111011011111,
24'b000000010001000001101011,
24'b001000110011111000101011,
24'b111111101101000011000010,
24'b110111111101000011100001,
24'b001010101011000010110111,
24'b111100010110111000011100,
24'b110001111000000000111100,
24'b010010101000000010000000,
24'b111111001110000010000010,
24'b110100011111111110100110,
24'b001001001001111110110111,
24'b110111010010111100011111,
24'b000111011100001001110000,
24'b000000101100111000100001,
24'b111101100011111111010100,
24'b111100111110000100110111,
24'b000010101110111100100010,
24'b111111101001000011001101,
24'b000110000101111011110010,
24'b110000100000000001100001,
24'b010010100000000000100000,
24'b110100101111000010000110,
24'b000001011101000000100011,
24'b111111101000110011101111,
24'b000010101111010011001100,
24'b000011010110110001010001,
24'b110110100100000111101010,
24'b000101010011111100100001,
24'b111101000010000011000010,
24'b001001010000111001011010,
24'b110110011001000111001000,
24'b111110111001000000000001,
24'b001010010111111010111110,
24'b110011111111000000101110,
24'b000111110001000110001000,
24'b000000001100110111000101,
24'b111101110001000101111100,
24'b111010100111000010101101,
24'b000101001111110110101101,
24'b001000011000000111000101,
24'b110100100000111011011100,
24'b000000001011001010101101,
24'b111110011100101101111110,
24'b001100001001001110110011,
24'b111100001110111111000011,
24'b110101001100110100101010,
24'b000100110101001001100000,
24'b000101010101000000110110,
24'b111101111111111110010010,
24'b000000001011111010010010,
24'b111100101100000011111101,
24'b000001111100000110000010,
24'b111101000010110111001110,
24'b000100010010000011001111,
24'b000101111111000000110111,
24'b110100001101000000010001,
24'b000000010101111100001100,
24'b000110110010000010101001,
24'b111110000101000101000011,
24'b000000110011111001110101,
24'b000000100101111001100010,
24'b111001011010010000010000,
24'b000010101111110100110101,
24'b000101100101000011101001,
24'b111110101000111100100011,
24'b111011010111000011011011,
24'b111111100010111111110000,
24'b000110111011111111000110,
24'b111010001110000000001100,
24'b111110111000000000010101,
24'b000101000010111101010100,
24'b000011010010000100001110,
24'b110100001111000000100101,
24'b000101111000111001010111,
24'b111110000101000110000011,
24'b000111001001111101000100,
24'b000000000101000010101000,
24'b110101011110111101101001,
24'b111101111100000011110110,
24'b010000000101110110110110,
24'b111000010001000101110000,
24'b111101111011001010010111,
24'b000011011000101110111001,
24'b111001000110000110000011,
24'b000100101001111111011101,
24'b000001111010001001010100,
24'b000011001101110011110010,
24'b111000100100000010100100,
24'b000001100110000011100111,
24'b111011111110000001010010,
24'b000110101101110111100111,
24'b000101101011001001101100,
24'b111010001100110111100001,
24'b110101101010001000100100,
24'b000010111111111110001100,
24'b010010011110110100010101,
24'b110011001010001011001100,
24'b111011101101000010111000,
24'b000110011111111101110101,
24'b111000000010110110000100,
24'b001001101011000110011100,
24'b000001000100000001100001,
24'b111011101111000100000001,
24'b110101011100111100000101,
24'b001111001100111001110101,
24'b111110100001000100001011,
24'b111001111010000010010011,
24'b000000011100000000111110,
24'b000110000001000001011010,
24'b111000101100111010010101,
24'b000010100001110111110111,
24'b000101100101010010001001,
24'b111001001000111110010101,
24'b111111001110110010101100,
24'b000100010110000110100001,
24'b000001110011000011000000,
24'b111011101011111100100011,
24'b111110011000111111011010,
24'b000001011101000100110001,
24'b000101001010111101001010,
24'b111101011010111110110100,
24'b111110000000111110001100,
24'b111100011111000001111101,
24'b000001100000000100111000,
24'b001011110101111011110011,
24'b111000011111000100000001,
24'b110101001101101110001101,
24'b001011001010010110001111,
24'b111111011001111000100001,
24'b000000000111000010101111,
24'b111111100000110111011110,
24'b111110011111000000111001,
24'b111101000000000111011111,
24'b000100000000111111010010,
24'b000010001011111011001101,
24'b111100101100000100111000,
24'b000100101100110111000110,
24'b110110000101000111000101,
24'b000110111101000001110101,
24'b111011001100111111000001,
24'b001011110010111010011101,
24'b111010111100000101000100,
24'b110101000010111101000010,
24'b000100001110111110110001,
24'b001000000001001101100010,
24'b000100011101101100001010,
24'b110000000010001010011100,
24'b000101110100000001010011,
24'b000011010011111000011010,
24'b111100111000001000100011,
24'b000011001101000001001001,
24'b111110000001110101111011,
24'b000100110001111110110110,
24'b110101000110001111100111,
24'b000000111101111000100110,
24'b001110011000111100011100,
24'b111000111110111011001001,
24'b111011001100000101111111,
24'b111111000111001101111011,
24'b111111101111101111001001,
24'b010000011101111001110110,
24'b101110110111001100001101,
24'b111101111111000011000011,
24'b001111010001111101101000,
24'b110101001011110111100001,
24'b111100000000000011001011,
24'b001011011010000011110000,
24'b111101101000000000010000,
24'b111011011010000000100111,
24'b111111000111111110000000,
24'b000000001111111001111010,
24'b000111000010000100010101,
24'b111101000001001000000101,
24'b111110110010111010100100,
24'b111000100000111011110100,
24'b001000100010000000001111,
24'b000110100111000100101001,
24'b110000001010111100010101,
24'b001010101101001000110101,
24'b111110000101110011000100,
24'b111100010000001011001010,
24'b000010111100101111001001,
24'b000001010011010010011101,
24'b111111010010000010110100,
24'b111111001100101010011001,
24'b111111001101001011011111,
24'b111011001100000111001101,
24'b001111101001110111010000,
24'b110011000010111110110110,
24'b111111110000000101000010,
24'b000010100111000001011000,
24'b000110101101111100000110,
24'b110100001001111011101011,
24'b001001101101000101011111,
24'b110111110101000110000110,
24'b000111100110110110100110,
24'b111110110001000010010011,
24'b110111111101111111001001,
24'b001000010000000001110001,
24'b111111101000111110110110,
24'b111101111000000110011100,
24'b000000100010111000111010,
24'b111001100111111011111001,
24'b001101100111000111111000,
24'b110111000101111101111011,
24'b000000101101000011100101,
24'b111100001100111011101101,
24'b001011000001111101100110,
24'b110111100001111111101011,
24'b000011101001000110011110,
24'b111001010100000010110001,
24'b000100001000110011111000,
24'b001100000111001000010011,
24'b101100111110111000011010,
24'b000110010010001011001001,
24'b000000111110111001000011,
24'b000101100001000011011010,
24'b111011000100111100100011,
24'b111101001100111100101000,
24'b000010101100000111100111,
24'b000000100110111111110101,
24'b111101101110111100010100,
24'b000101101110000001001000,
24'b111111000111111010001110,
24'b110100110000001010011001,
24'b001001101100111011011110,
24'b111111110001111111111110,
24'b000010010111000001001111,
24'b111110111000110100001111,
24'b110100110101010100110000,
24'b000101111111110111011111,
24'b001101110001110110000010,
24'b110100111011001001000001,
24'b111001011110000010011011,
24'b000101111010111101011100,
24'b000011100111111101110000,
24'b111111101011111100101010,
24'b111010111000001001110010,
24'b000000010011111100110110,
24'b000110111001111010000000,
24'b110110110001000101100100,
24'b000111010100111100001010,
24'b111100101010000101000011,
24'b000010000001000010001100,
24'b111011100000110001101111,
24'b000011110101001011001110,
24'b000011110001000100000110,
24'b110110011110110111101010,
24'b000101000011000001000001,
24'b000000110001111111011010,
24'b000011101110000101010101,
24'b111000111011111010111110,
24'b111011101101001000001011,
24'b001100111100110001110110,
24'b111110010100000011001101,
24'b110111101000001111011010,
24'b111110110110110011110011,
24'b001001101011000000011100,
24'b111110010101111000111010,
24'b111010011010001100000110,
24'b000011111100000001100000,
24'b111001000011111011001110,
24'b001101101011110111000111,
24'b110100100001001000000011,
24'b000101110001000011110100,
24'b111011011111111111100101,
24'b111110101011111001101100,
24'b001011011011000000111010,
24'b110101110011111111011010,
24'b000001011101001001000000,
24'b000000000000111001010010,
24'b000000011101111100100010,
24'b000000110100000101110101,
24'b000110111110111101001100,
24'b110100010000000000011000,
24'b111011001110000000111101,
24'b010011111001000011000000,
24'b110011101011111000110011,
24'b000011101100000001010011,
24'b111010100110000011111111,
24'b000011010110000011111101,
24'b111100010101110100101110,
24'b001010001110001000000010,
24'b111101110110111001100011,
24'b110100000111001001000001,
24'b000100101110111000010011,
24'b000101111101000111001010,
24'b111111110111111001000011,
24'b000010000111111110010110,
24'b101111110001000111010100,
24'b001100001110111111100101,
24'b000100110010111111000111,
24'b111000110000111001101000,
24'b000000110000000001110110,
24'b000000001101000110010010,
24'b111111101111111111010111,
24'b000010011010111101100011,
24'b111110001011111011101110,
24'b111100100000000010001100,
24'b001010011111000100100000,
24'b110101100100111100010010,
24'b000011110111000110001101,
24'b111011110110111000101100,
24'b000111100010111100010101,
24'b000000011000000011010110,
24'b111010010001001011000000,
24'b111000101101111100001111,
24'b010001101110110001000101,
24'b110111011000001010010011,
24'b111110001100111101000100,
24'b111111101010001011100010,
24'b000101101100110101010001,
24'b111001101001000010111111,
24'b000101000010111001110100,
24'b111010110001000000011100,
24'b000101101111001100110101,
24'b111011011010111010110000,
24'b000110011000111101110011,
24'b110100110111110101000011,
24'b000111000010001000101000,
24'b000100011110001100010001,
24'b111000100111110100100000,
24'b000100001101000000000101,
24'b111010111001111011101110,
24'b000011101111000011101011,
24'b111110100111000110111010,
24'b001000000111111001110011,
24'b110010010011000010010111,
24'b001001100100111101100100,
24'b111011000010111001010001,
24'b111100011001001011100001,
24'b010010011000000001000001,
24'b101110110110111010001100,
24'b000000111111111100100000,
24'b000001011000000100010111,
24'b000101110101000000001011,
24'b111100010100000000010010,
24'b000010001111000010011010,
24'b111100110011111101001101,
24'b111010011011111001100100,
24'b000111100000000111100001,
24'b001000011011000011010100,
24'b110000111001111010111100,
24'b000011110101111100011100,
24'b000010010000000110011001,
24'b000000100111000000111100,
24'b111101111001110010101011,
24'b000011000100010011000101,
24'b111111110101110110100001,
24'b111000000101111111001111,
24'b001001001011111101111100,
24'b111010001001000010000110,
24'b001010001011001010010111,
24'b110110000110110001110100,
24'b111000111000000000110011,
24'b010100001011000011001001,
24'b110010011101010000101000,
24'b000110000011100011000010,
24'b110110100111000110101001,
24'b000100010111010011000110,
24'b001101011100110110110100,
24'b110010110110110110000110,
24'b110001101110000001011000,
24'b011111001100000111001000,
24'b101110000110001011000000,
24'b000010001010101011111101,
24'b111110010000111110010000,
24'b000100001000010010101010,
24'b111101000001110101101110,
24'b000001000111111101101111,
24'b000010111000000101111101,
24'b111100000101111100000111,
24'b111110110011111011000111,
24'b000011001111001101001111,
24'b000000100110111011000010,
24'b111011000010110010101111,
24'b001001000101001101100101,
24'b110111000010000101101001,
24'b000100110100110011010001,
24'b111001100001111111010011,
24'b000110010111000111111101,
24'b000100101100111101000111,
24'b111101011111000010010101,
24'b101101111000111110000011,
24'b010001111111111100101010,
24'b000011100100111101011110,
24'b111010000100001100101111,
24'b111011000001111100000100,
24'b000011100111110111011001,
24'b111011100010000011001101,
24'b001011010010000101011110,
24'b111100100000110110110000,
24'b111010110111001110100110,
24'b111100001100111000011001,
24'b000111001001110110011110,
24'b000111010111000110011000,
24'b101111110010001000010100,
24'b001001011001111101000011,
24'b000000100000111001101001,
24'b111100110111111111000001,
24'b111101111010000010011011,
24'b000100101100001000011011,
24'b000000011000110111101101,
24'b111111011000000010101000,
24'b111010110000111001000001,
24'b000100110011000110110011,
24'b111101000011000100000010,
24'b000100111010111001111101,
24'b000001100100111111001111,
24'b110011001101111110010001,
24'b001100010111001010000101,
24'b111100000100110110010101,
24'b111011111010000011101010,
24'b000111010011111110000101,
24'b000100100010000011101110,
24'b101101101011111100101100,
24'b000111001111111101101110,
24'b001010111011001001101000,
24'b111010111000110111111011,
24'b111001100101111011111001,
24'b000001001110001010001110,
24'b000110000111111101101010,
24'b111010010000111011000111,
24'b000011011011000100111100,
24'b000000011010111001110110,
24'b111111010111000100101010,
24'b111011011000000010101000,
24'b000100000001111110111111,
24'b000000011000111000011100,
24'b000001010100000011100000,
24'b111110000110000101110111,
24'b000000000000111011000011,
24'b111110001011000101001001,
24'b111100101000110110011010,
24'b001100100010000100001000,
24'b111011101000000001011011,
24'b111001111000000111000101,
24'b111011111010110000111010,
24'b001011101110001100100111,
24'b111101011110111010110001,
24'b000000100101111000100101,
24'b111000110110001110011101,
24'b000111010101111110001011,
24'b111000011110110111000000,
24'b000100011100000000100010,
24'b001000000111000100010001,
24'b111000010001000001100100,
24'b111010110110000010100110,
24'b000010011101110111011101,
24'b000010100000000000100010,
24'b000110011101000101110010,
24'b000000100000111011110110,
24'b101111101000001000110010,
24'b111111110110110010001011,
24'b010011001100000111011001,
24'b111110100110000001100000,
24'b110111110011111011100010,
24'b110100010100000011001000,
24'b001001110001000000010001,
24'b001011100010000000000001,
24'b111001011111111101010010,
24'b111011110101111101011100,
24'b111100001011001010011010,
24'b111101010111110111101101,
24'b010011001100000011010100,
24'b111001100010111100001111,
24'b110111101111000011000100,
24'b110111101110000001100100,
24'b001101100000111010011001,
24'b001100011010000110100001,
24'b101011001010111100010111,
24'b000100100110000010100001,
24'b111101101010111010000100,
24'b000110000000000100101100,
24'b000110000110111110011101,
24'b110101110010000111101001,
24'b111100100011111000111101,
24'b000111001101110110000100,
24'b000001101011001011100100,
24'b111001111000001001110000,
24'b001001100110110001101000,
24'b110110110000111110010110,
24'b111000001100000010010101,
24'b010110100101001100000010,
24'b110100111111110010000101,
24'b110111110100000001001101,
24'b001010011110000111110001,
24'b111101110000000000100110,
24'b111010000011110000011101,
24'b001011010101001001111010,
24'b110111110100001000011100,
24'b000000111000111010100110,
24'b111110111011111000011001,
24'b000011011111000010010000,
24'b000010111101000010111100,
24'b110011100010000011110100,
24'b001111100110000001011111,
24'b110011111010110111001110,
24'b000100000111111010110110,
24'b000001101100001101000111,
24'b000100011001111111101111,
24'b101111001100111101111111,
24'b010000101001111010111000,
24'b111110010101111101000011,
24'b111000111101001001110111,
24'b111110111001111011010110,
24'b001000011110001000000010,
24'b111101111001110100011111,
24'b111110110000111101101010,
24'b110110100101001010110101,
24'b001100111010111100101100,
24'b000001100000000000000001,
24'b110111010100000001101100,
24'b111101001010111000101101,
24'b001001010111111111110011,
24'b111101111000001001001000,
24'b111111100010000011010010,
24'b111100010010110100101111,
24'b000011001001111110011100,
24'b111011011100000010100110,
24'b001011010001001000110100,
24'b111011101110111111100000,
24'b110001011011110101011111,
24'b001111011011111101010111,
24'b000001010101001101110010,
24'b111010111101111010110101,
24'b111011111010111111101111,
24'b000011001011111011011101,
24'b000100010001001000100010,
24'b111011100100110100110110,
24'b000010000010001001011100,
24'b111110111100111011000111,
24'b111111110100001011000101,
24'b111101000110101100101001,
24'b000101010001001011110110,
24'b000100010010111101000001,
24'b110010111010000100100100,
24'b000101110001111110000100,
24'b000011010110111101010010,
24'b111110011000111111001111,
24'b111110011010111111111001,
24'b000100100010000100010001,
24'b110111011011000001011101,
24'b000000111101111110101100,
24'b001101000101111000010110,
24'b110110011011111101001111,
24'b111111000001010101010111,
24'b111000011010101111011011,
24'b010010000101000110111111,
24'b110111100111111000011110,
24'b000011100011111010111110,
24'b101110111110010011010001,
24'b001111001001111000110010,
24'b000110111111111001011111,
24'b110110001001000001001010,
24'b111010010001000001000101,
24'b000101001010000010111110,
24'b000001100001111101101111,
24'b001001001010000111100111,
24'b110000111010110010111100,
24'b000011110010000010001000,
24'b111100110011000110110101,
24'b001101100101111110010111,
24'b110111000011111111110000,
24'b000000011000000000110111,
24'b111011000010111001100011,
24'b000100101100111111011101,
24'b000100110101001100010101,
24'b111100001111111100001011,
24'b111101001001111000100001,
24'b000001110101111111101110,
24'b111101110001001001011111,
24'b000100001000111000010100,
24'b000011101010000010010010,
24'b110100000100000011001110,
24'b001010000111111111110100,
24'b111010010101110100110110,
24'b000010000000001001100001,
24'b000010101111000001101110,
24'b111100010111000000110001,
24'b000000010011111010001010,
24'b000010110010111111001101,
24'b111011100101000001100001,
24'b000001001110000100000010,
24'b000100011100000010010111,
24'b111101010101110110010000,
24'b111110101110000100100111,
24'b111101000111000001101110,
24'b000101001000111011110101,
24'b000001001010000011110111,
24'b111011100011000010001111,
24'b000000111010111110000111,
24'b000101010000110110011110,
24'b110100010000001001110110,
24'b001000011110000001000111,
24'b000100111000111111010011,
24'b110111000010111100101000,
24'b000001110110111110001010,
24'b000010001000000000110110,
24'b111100010010000101110100,
24'b000010010111000001000111,
24'b000100000111110100111111,
24'b000001101010000110000001,
24'b110000110011000001111101,
24'b000101011110111111000010,
24'b001100000110111110000111,
24'b111010100000000000001101,
24'b000001101110000110000010,
24'b101110000011110011110101,
24'b010001110111001010011000,
24'b111110001111111101100101,
24'b000010011101111101001110,
24'b111000101100000011000000,
24'b000011110001111111111111,
24'b110111000101111101110001,
24'b001001010111111101101101,
24'b000110011000001000110010,
24'b111010011101111001001011,
24'b110110001000111111000011,
24'b000100100011000111000000,
24'b000100001100110111110111,
24'b000011010000000001010010,
24'b000010001101000111100010,
24'b110001111110111000101010,
24'b111101101010000101101001,
24'b010010000010110011111101,
24'b111110010111001101111110,
24'b110110000011111101110001,
24'b111101101011110100111000,
24'b000101101100010000001000,
24'b000101101001110100111010,
24'b110110001111111101001110,
24'b000110000111001100111000,
24'b000000101100110111110101,
24'b110011101011111110110110,
24'b010000110000000010010001,
24'b111011000010000000111100,
24'b111001010001000000001111,
24'b000010010011111100110111,
24'b000111100110111101001101,
24'b111010110011001101100010,
24'b111101101000110111011110,
24'b111110000001111000001000,
24'b001000101100000111100101,
24'b111110010101000001110110,
24'b111010000011000101110010,
24'b000010110111110100001110,
24'b111100011011111101100011,
24'b001001111100000111001001,
24'b111000101011000100101101,
24'b000001101100000000011110,
24'b111100101011110001001101,
24'b000011001110000110101001,
24'b000011110111000111000000,
24'b110011001101111101100000,
24'b010011101101111011111000,
24'b101111111001000010001111,
24'b000100100011111101100101,
24'b111001000010000101101001,
24'b010011011000111000010101,
24'b110011111010001000010100,
24'b111000111100111011000000,
24'b000110000111000000000101,
24'b000111110100000001011110,
24'b110110111111000000100011,
24'b000000111110110101100010,
24'b000010111010010110101101,
24'b111100011101110001011000,
24'b000100010000111000111110,
24'b111101011110000111011100,
24'b111011101110000110001110,
24'b001011101000111111110000,
24'b110101010110110001101111,
24'b000100100011001001011111,
24'b111011111111000011011101,
24'b000100110010111011011101,
24'b000000001010111100010100,
24'b111111100011001011110110,
24'b111001010011110100010010,
24'b000100110011000011001110,
24'b000111110001000000111111,
24'b110100010000000001100011,
24'b000010111110000000101000,
24'b000010000100111001001111,
24'b000011011111000111110001,
24'b111001110010111101111000,
24'b111111000111110111011011,
24'b000010111101001110011000,
24'b000101110100111010111101,
24'b111100100000111101111011,
24'b110001100010111001011100,
24'b010010100000000101100001,
24'b111101001010001010000001,
24'b111011000011111110110110,
24'b000010100010100101101010,
24'b111001001011010110010001,
24'b001000000010000011110110,
24'b000100110010111011111111,
24'b110010011000110101100100,
24'b001000110010000101100000,
24'b111100100000000100001110,
24'b000000010111111110111110,
24'b000111001001000001010100,
24'b110101010011111000001110,
24'b000010111010000000011011,
24'b000011110111001111100101,
24'b000000101101110001110010,
24'b111001111111111101111011,
24'b000001110101000110010100,
24'b000001110110000010101100,
24'b000100000110000000010111,
24'b110111100101110010111101,
24'b000011100001000110101111,
24'b000000101000001011111011,
24'b111100110101110011111000,
24'b001100110010000011010000,
24'b101110110100110111110100,
24'b000010001101001000001110,
24'b001100001101001001100101,
24'b111011100111110000010010,
24'b111000010001000000001111,
24'b000010100011001010010110,
24'b000110001101111000010011,
24'b111110011010000000101011,
24'b111010101010001001101011,
24'b000010110100110011011000,
24'b000000011110000010010010,
24'b000001111010000000110000,
24'b111100001001000111101001,
24'b000100110010111000100110,
24'b111000110011000101111100,
24'b000101011100110000110110,
24'b111111101000001100110110,
24'b000010000100000010001111,
24'b111010110000000000000110,
24'b111110011101110101101101,
24'b000111110101000010010001,
24'b111110111000000100110001,
24'b111000101001000011000010,
24'b000111101011111110110111,
24'b111001100100110100100110,
24'b000101011001001110100010,
24'b111111111110110000110000,
24'b111010001011010001001111,
24'b000111011100111010001110,
24'b111001011111111001111111,
24'b000101100011111101101010,
24'b111001101100001100100011,
24'b000110010001111001011101,
24'b000001001101111110100011,
24'b110101000010000001011010,
24'b001001110010000000100101,
24'b111111001000111110100001,
24'b111110010101000000101100,
24'b111101010010111110101100,
24'b000110100011000111110100,
24'b110111111111110111101110,
24'b000110010000111011011110,
24'b111111010000001000100001,
24'b111101111011000011110111,
24'b111110010010111100010010,
24'b000011010100110101000111,
24'b000100010101000100000111,
24'b110110111100010011100011,
24'b111110111111110001000100,
24'b001010101101110000001000,
24'b111011110010010111001100,
24'b111110111110000010000111,
24'b111000011010101101001101,
24'b001001000001001000101111,
24'b000000111000000110100110,
24'b000001111101110101000011,
24'b110101010010000100011000,
24'b000011001101001000111001,
24'b000011000010110001000001,
24'b000110101010000100111101,
24'b110111001000000100011101,
24'b000000010000000000101100,
24'b111111111100111000110011,
24'b111111000111000100101000,
24'b001000001000000001101100,
24'b111111010100110110111000,
24'b110110000010001100101110,
24'b111100111101111000111101,
24'b001111100010000010100000,
24'b111100001111111101101110,
24'b111100000000111000010001,
24'b111100011101010001011011,
24'b000010111000111010011101,
24'b000001001010110111010111,
24'b000100110111000011101010,
24'b111100100101111111010111};