logic pilot [0:71] = {
1,
0,
0,
1,
1,
1,
0,
1,
1,
0,
1,
0,
1,
0,
0,
1,
0,
0,
0,
0,
1,
1,
0,
1,
1,
1,
0,
1,
1,
0,
0,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
0,
0,
0,
1,
1,
1,
1,
0,
1,
0,
1,
1,
1,
1,
0,
1,
1,
1,
0,
0,
1,
1,
1,
1,
1,
0,
0,
0,
0};