logic [23:0] rom_freq_pr [0:6143] = {
24'b111000011001001000110101,
24'b000111101001111010100000,
24'b111101000100111000100000,
24'b000101110001001011100110,
24'b111101100010110011001011,
24'b111000010100001111100101,
24'b001000010001110111000111,
24'b111011100011111110111011,
24'b000100010001000010010011,
24'b000001100000111111100010,
24'b111000100111111110110111,
24'b000001011001000011011110,
24'b000001111100000010011011,
24'b000101111101110011001011,
24'b111100001100001010101000,
24'b110011110111111110010100,
24'b010000101000000010100100,
24'b111011100000111011001111,
24'b111101000000111101110101,
24'b111100110101000011000101,
24'b001100100100001100110011,
24'b110001001111100101110101,
24'b001001100111010000011110,
24'b111100101100000011101001,
24'b111111101101111000111100,
24'b000001111100111100011011,
24'b111111100110000100011000,
24'b111010000001000011100011,
24'b001100110000111111101000,
24'b110011011011110101101000,
24'b000100100000001010100001,
24'b000011100111111111111001,
24'b111010101111111001110000,
24'b000011010101111111001101,
24'b111111011000001101000000,
24'b111100111110110111000111,
24'b111111110101110101101111,
24'b001010001101001101101000,
24'b111001110110000010011011,
24'b110101010101111010000000,
24'b000111001011111011110101,
24'b001100000010000010001011,
24'b110110011001000011100101,
24'b111101001110000110011011,
24'b111011111000110001110110,
24'b000101100000000100000101,
24'b001111001101000101010000,
24'b101011100111111100000100,
24'b000001011011000011110100,
24'b000110011101111011100010,
24'b111111110011111101110110,
24'b111100001011001001101011,
24'b001010101011110110011111,
24'b110001100000000100011001,
24'b000011000010111111011111,
24'b000110000101000000111100,
24'b111110000111111101000001,
24'b000011010011000001110000,
24'b110110011111111111001001,
24'b000000100011000101101001,
24'b001101110110110111001001,
24'b110111100001000011100111,
24'b110011101110000010101111,
24'b010101000110111011111111,
24'b110111011000000011011111,
24'b111101001001111101010010,
24'b111110101100000011001001,
24'b000100101010110111010010,
24'b111111000010001101100111,
24'b000011111010110111100010,
24'b111011100100111111101110,
24'b111010010100000000101000,
24'b000010110011000101101010,
24'b001011000101110110000010,
24'b111000101100001000010010,
24'b000001000100111100101011,
24'b110110110001000010100010,
24'b000001101001111100000011,
24'b010000100101111101001111,
24'b111001011000001001001010,
24'b111001001001000000011110,
24'b111000001001110111001001,
24'b001111010111111010111101,
24'b111100110000010001100000,
24'b000011100100111010011100,
24'b111001111000111001101110,
24'b111001110010111110001001,
24'b001001101000001011001011,
24'b111100110001110110011010,
24'b000011100001000111001001,
24'b000100001000111011000000,
24'b110001010110111110001010,
24'b000100100100000110110100,
24'b000010101001111111111111,
24'b001001101100110001010001,
24'b110110010001010001000110,
24'b111110011100000001011011,
24'b111100000110110010111101,
24'b001010001101111111010011,
24'b111011100100001010001001,
24'b000101111101000000101101,
24'b110111101110111101110110,
24'b111111000111110111001011,
24'b000011010000000011101001,
24'b000000111000000111001101,
24'b000011110100111110110100,
24'b111011110010111011011000,
24'b111100100111000001111111,
24'b000001110101111010001010,
24'b000001011011000110010001,
24'b000010111110000011010010,
24'b111101111001000001110000,
24'b111111110011101110101101,
24'b111010101011001110001100,
24'b000101010101111100111101,
24'b000000100001000011010110,
24'b000000100011111111111100,
24'b111111100010110110001011,
24'b111011100000001000111011,
24'b000100111101111101100000,
24'b111000110001000001010100,
24'b001011010111111111011000,
24'b111100010010000010010010,
24'b111100101000111001111110,
24'b111011011000000001010101,
24'b001011100101000101001111,
24'b110101011000111100111011,
24'b001010011000000010010010,
24'b111000111101111010000100,
24'b000100001011000111010111,
24'b111000110000110011111101,
24'b000001111101001101111011,
24'b000100000101111110000111,
24'b001010010011111100101010,
24'b101100011110111010110001,
24'b000101000000111101101000,
24'b000000001101010000100000,
24'b000011100000111100001011,
24'b001101110010111000000101,
24'b100111000101111011000000,
24'b000110111101000010011000,
24'b000001111001010010100001,
24'b000101011011110011010011,
24'b000000110100111100110111,
24'b111001010011111010101111,
24'b000000100110000111101101,
24'b111000111011001000100111,
24'b001110001110110111010110,
24'b000001101100000000001100,
24'b110110000101110110111111,
24'b111100011010001001010101,
24'b000000100001001100111010,
24'b010010011011101000111000,
24'b110011100100001001111011,
24'b110110010101000100000000,
24'b001000100111110111101100,
24'b001000101100000011011101,
24'b110101111011000110000010,
24'b000010000000111000001110,
24'b110101101100000010111111,
24'b010101111010111101000110,
24'b110101100010000100101100,
24'b111010010100111011110110,
24'b000011001110000100111100,
24'b111111110111111010111101,
24'b000100100100000101011010,
24'b111110100000110111000000,
24'b000010011101000101011110,
24'b110100001001000011011011,
24'b000000010110000011010010,
24'b010011111110101111000101,
24'b111000101101001010111011,
24'b101111010001000001100110,
24'b001101000001000010010101,
24'b111111101010110111111001,
24'b111101111011000010011010,
24'b000110000000000001101000,
24'b110100111101000000011010,
24'b001011101000000000011010,
24'b111000100010111011101011,
24'b111000101011000111011001,
24'b010000111100111001100001,
24'b111100110001000000000110,
24'b111010001011000100011101,
24'b111011001011111101111110,
24'b000100101101000001011111,
24'b000010100011111000100101,
24'b000100001011001001101011,
24'b000001100101111110100010,
24'b101100110000111001010011,
24'b000100110010000000001111,
24'b010100100000001010100101,
24'b110100100000111111110001,
24'b111110001101101101100111,
24'b111010101111001010011010,
24'b000011101011000101011001,
24'b000110001010000101001011,
24'b111001100010110101010111,
24'b001011100111110010100101,
24'b101110001111010100110101,
24'b000101111111111111001101,
24'b000111000010000011101111,
24'b110110011110101010111111,
24'b001100111001000111111011,
24'b110110100101001000110101,
24'b111110110110000100000010,
24'b000000000100110011110011,
24'b000010100100111101011010,
24'b000000111101001010101101,
24'b001011110111111001011000,
24'b100110000010000100110010,
24'b001001010111111110111001,
24'b001000111101111011110100,
24'b111100001110000100011001,
24'b000100010010111011001101,
24'b110100000011000011100101,
24'b000010101000000100100000,
24'b000101010001111000101111,
24'b000001100001000010101001,
24'b000001011110111010011011,
24'b110100001110001011100000,
24'b000111100111110110101011,
24'b000000000111000110110111,
24'b000001011111111011111011,
24'b111101100011111011011001,
24'b111110001100000100110101,
24'b000111001011000100100001,
24'b111000001001111110100101,
24'b000000011010111001010110,
24'b000000011000111101111011,
24'b001101111011001011001100,
24'b101110100000111011011111,
24'b000000010001000001101011,
24'b001000110011111000101011,
24'b111111101101000011000010,
24'b110111111101000011100001,
24'b001010101011000010110111,
24'b111100010110111000011100,
24'b110001111000000000111100,
24'b010010101000000010000000,
24'b111111001110000010000010,
24'b110100011111111110100110,
24'b001001001001111110110111,
24'b110111010010111100011111,
24'b000111011100001001110000,
24'b000000101100111000100001,
24'b111101100011111111010100,
24'b111100111110000100110111,
24'b000010101110111100100010,
24'b111111101001000011001101,
24'b000110000101111011110010,
24'b110000100000000001100001,
24'b010010100000000000100000,
24'b110100101111000010000110,
24'b000001011101000000100011,
24'b111111101000110011101111,
24'b000010101111010011001100,
24'b000011010110110001010001,
24'b110110100100000111101010,
24'b000101010011111100100001,
24'b111101000010000011000010,
24'b001001010000111001011010,
24'b110110011001000111001000,
24'b111110111001000000000001,
24'b001010010111111010111110,
24'b110011111111000000101110,
24'b000111110001000110001000,
24'b000000001100110111000101,
24'b111101110001000101111100,
24'b111010100111000010101101,
24'b000101001111110110101101,
24'b001000011000000111000101,
24'b110100100000111011011100,
24'b000000001011001010101101,
24'b111110011100101101111110,
24'b001100001001001110110011,
24'b111100001110111111000011,
24'b110101001100110100101010,
24'b000100110101001001100000,
24'b000101010101000000110110,
24'b111101111111111110010010,
24'b000000001011111010010010,
24'b111100101100000011111101,
24'b000001111100000110000010,
24'b111101000010110111001110,
24'b000100010010000011001111,
24'b000101111111000000110111,
24'b110100001101000000010001,
24'b000000010101111100001100,
24'b000110110010000010101001,
24'b111110000101000101000011,
24'b000000110011111001110101,
24'b000000100101111001100010,
24'b111001011010010000010000,
24'b000010101111110100110101,
24'b000101100101000011101001,
24'b111110101000111100100011,
24'b111011010111000011011011,
24'b111111100010111111110000,
24'b000110111011111111000110,
24'b111010001110000000001100,
24'b111110111000000000010101,
24'b000101000010111101010100,
24'b000011010010000100001110,
24'b110100001111000000100101,
24'b000101111000111001010111,
24'b111110000101000110000011,
24'b000111001001111101000100,
24'b000000000101000010101000,
24'b110101011110111101101001,
24'b111101111100000011110110,
24'b010000000101110110110110,
24'b111000010001000101110000,
24'b111101111011001010010111,
24'b000011011000101110111001,
24'b111001000110000110000011,
24'b000100101001111111011101,
24'b000001111010001001010100,
24'b000011001101110011110010,
24'b111000100100000010100100,
24'b000001100110000011100111,
24'b111011111110000001010010,
24'b000110101101110111100111,
24'b000101101011001001101100,
24'b111010001100110111100001,
24'b110101101010001000100100,
24'b000010111111111110001100,
24'b010010011110110100010101,
24'b110011001010001011001100,
24'b111011101101000010111000,
24'b000110011111111101110101,
24'b111000000010110110000100,
24'b001001101011000110011100,
24'b000001000100000001100001,
24'b111011101111000100000001,
24'b110101011100111100000101,
24'b001111001100111001110101,
24'b111110100001000100001011,
24'b111001111010000010010011,
24'b000000011100000000111110,
24'b000110000001000001011010,
24'b111000101100111010010101,
24'b000010100001110111110111,
24'b000101100101010010001001,
24'b111001001000111110010101,
24'b111111001110110010101100,
24'b000100010110000110100001,
24'b000001110011000011000000,
24'b111011101011111100100011,
24'b111110011000111111011010,
24'b000001011101000100110001,
24'b000101001010111101001010,
24'b111101011010111110110100,
24'b111110000000111110001100,
24'b111100011111000001111101,
24'b000001100000000100111000,
24'b001011110101111011110011,
24'b111000011111000100000001,
24'b110101001101101110001101,
24'b001011001010010110001111,
24'b111111011001111000100001,
24'b000000000111000010101111,
24'b111111100000110111011110,
24'b111110011111000000111001,
24'b111101000000000111011111,
24'b000100000000111111010010,
24'b000010001011111011001101,
24'b111100101100000100111000,
24'b000100101100110111000110,
24'b110110000101000111000101,
24'b000110111101000001110101,
24'b111011001100111111000001,
24'b001011110010111010011101,
24'b111010111100000101000100,
24'b110101000010111101000010,
24'b000100001110111110110001,
24'b001000000001001101100010,
24'b000100011101101100001010,
24'b110000000010001010011100,
24'b000101110100000001010011,
24'b000011010011111000011010,
24'b111100111000001000100011,
24'b000011001101000001001001,
24'b111110000001110101111011,
24'b000100110001111110110110,
24'b110101000110001111100111,
24'b000000111101111000100110,
24'b001110011000111100011100,
24'b111000111110111011001001,
24'b111011001100000101111111,
24'b111111000111001101111011,
24'b111111101111101111001001,
24'b010000011101111001110110,
24'b101110110111001100001101,
24'b111101111111000011000011,
24'b001111010001111101101000,
24'b110101001011110111100001,
24'b111100000000000011001011,
24'b001011011010000011110000,
24'b111101101000000000010000,
24'b111011011010000000100111,
24'b111111000111111110000000,
24'b000000001111111001111010,
24'b000111000010000100010101,
24'b111101000001001000000101,
24'b111110110010111010100100,
24'b111000100000111011110100,
24'b001000100010000000001111,
24'b000110100111000100101001,
24'b110000001010111100010101,
24'b001010101101001000110101,
24'b111110000101110011000100,
24'b111100010000001011001010,
24'b000010111100101111001001,
24'b000001010011010010011101,
24'b111111010010000010110100,
24'b111111001100101010011001,
24'b111111001101001011011111,
24'b111011001100000111001101,
24'b001111101001110111010000,
24'b110011000010111110110110,
24'b111111110000000101000010,
24'b000010100111000001011000,
24'b000110101101111100000110,
24'b110100001001111011101011,
24'b001001101101000101011111,
24'b110111110101000110000110,
24'b000111100110110110100110,
24'b111110110001000010010011,
24'b110111111101111111001001,
24'b001000010000000001110001,
24'b111111101000111110110110,
24'b111101111000000110011100,
24'b000000100010111000111010,
24'b111001100111111011111001,
24'b001101100111000111111000,
24'b110111000101111101111011,
24'b000000101101000011100101,
24'b111100001100111011101101,
24'b001011000001111101100110,
24'b110111100001111111101011,
24'b000011101001000110011110,
24'b111001010100000010110001,
24'b000100001000110011111000,
24'b001100000111001000010011,
24'b101100111110111000011010,
24'b000110010010001011001001,
24'b000000111110111001000011,
24'b000101100001000011011010,
24'b111011000100111100100011,
24'b111101001100111100101000,
24'b000010101100000111100111,
24'b000000100110111111110101,
24'b111101101110111100010100,
24'b000101101110000001001000,
24'b111111000111111010001110,
24'b110100110000001010011001,
24'b001001101100111011011110,
24'b111111110001111111111110,
24'b000010010111000001001111,
24'b111110111000110100001111,
24'b110100110101010100110000,
24'b000101111111110111011111,
24'b001101110001110110000010,
24'b110100111011001001000001,
24'b111001011110000010011011,
24'b000101111010111101011100,
24'b000011100111111101110000,
24'b111111101011111100101010,
24'b111010111000001001110010,
24'b000000010011111100110110,
24'b000110111001111010000000,
24'b110110110001000101100100,
24'b000111010100111100001010,
24'b111100101010000101000011,
24'b000010000001000010001100,
24'b111011100000110001101111,
24'b000011110101001011001110,
24'b000011110001000100000110,
24'b110110011110110111101010,
24'b000101000011000001000001,
24'b000000110001111111011010,
24'b000011101110000101010101,
24'b111000111011111010111110,
24'b111011101101001000001011,
24'b001100111100110001110110,
24'b111110010100000011001101,
24'b110111101000001111011010,
24'b111110110110110011110011,
24'b001001101011000000011100,
24'b111110010101111000111010,
24'b111010011010001100000110,
24'b000011111100000001100000,
24'b111001000011111011001110,
24'b001101101011110111000111,
24'b110100100001001000000011,
24'b000101110001000011110100,
24'b111011011111111111100101,
24'b111110101011111001101100,
24'b001011011011000000111010,
24'b110101110011111111011010,
24'b000001011101001001000000,
24'b000000000000111001010010,
24'b000000011101111100100010,
24'b000000110100000101110101,
24'b000110111110111101001100,
24'b110100010000000000011000,
24'b111011001110000000111101,
24'b010011111001000011000000,
24'b110011101011111000110011,
24'b000011101100000001010011,
24'b111010100110000011111111,
24'b000011010110000011111101,
24'b111100010101110100101110,
24'b001010001110001000000010,
24'b111101110110111001100011,
24'b110100000111001001000001,
24'b000100101110111000010011,
24'b000101111101000111001010,
24'b111111110111111001000011,
24'b000010000111111110010110,
24'b101111110001000111010100,
24'b001100001110111111100101,
24'b000100110010111111000111,
24'b111000110000111001101000,
24'b000000110000000001110110,
24'b000000001101000110010010,
24'b111111101111111111010111,
24'b000010011010111101100011,
24'b111110001011111011101110,
24'b111100100000000010001100,
24'b001010011111000100100000,
24'b110101100100111100010010,
24'b000011110111000110001101,
24'b111011110110111000101100,
24'b000111100010111100010101,
24'b000000011000000011010110,
24'b111010010001001011000000,
24'b111000101101111100001111,
24'b010001101110110001000101,
24'b110111011000001010010011,
24'b111110001100111101000100,
24'b111111101010001011100010,
24'b000101101100110101010001,
24'b111001101001000010111111,
24'b000101000010111001110100,
24'b111010110001000000011100,
24'b000101101111001100110101,
24'b111011011010111010110000,
24'b000110011000111101110011,
24'b110100110111110101000011,
24'b000111000010001000101000,
24'b000100011110001100010001,
24'b111000100111110100100000,
24'b000100001101000000000101,
24'b111010111001111011101110,
24'b000011101111000011101011,
24'b111110100111000110111010,
24'b001000000111111001110011,
24'b110010010011000010010111,
24'b001001100100111101100100,
24'b111011000010111001010001,
24'b111100011001001011100001,
24'b010010011000000001000001,
24'b101110110110111010001100,
24'b000000111111111100100000,
24'b000001011000000100010111,
24'b000101110101000000001011,
24'b111100010100000000010010,
24'b000010001111000010011010,
24'b111100110011111101001101,
24'b111010011011111001100100,
24'b000111100000000111100001,
24'b001000011011000011010100,
24'b110000111001111010111100,
24'b000011110101111100011100,
24'b000010010000000110011001,
24'b000000100111000000111100,
24'b111101111001110010101011,
24'b000011000100010011000101,
24'b111111110101110110100001,
24'b111000000101111111001111,
24'b001001001011111101111100,
24'b111010001001000010000110,
24'b001010001011001010010111,
24'b110110000110110001110100,
24'b111000111000000000110011,
24'b010100001011000011001001,
24'b110010011101010000101000,
24'b000110000011100011000010,
24'b110110100111000110101001,
24'b000100010111010011000110,
24'b001101011100110110110100,
24'b110010110110110110000110,
24'b110001101110000001011000,
24'b011111001100000111001000,
24'b101110000110001011000000,
24'b000010001010101011111101,
24'b111110010000111110010000,
24'b000100001000010010101010,
24'b111101000001110101101110,
24'b000001000111111101101111,
24'b000010111000000101111101,
24'b111100000101111100000111,
24'b111110110011111011000111,
24'b000011001111001101001111,
24'b000000100110111011000010,
24'b111011000010110010101111,
24'b001001000101001101100101,
24'b110111000010000101101001,
24'b000100110100110011010001,
24'b111001100001111111010011,
24'b000110010111000111111101,
24'b000100101100111101000111,
24'b111101011111000010010101,
24'b101101111000111110000011,
24'b010001111111111100101010,
24'b000011100100111101011110,
24'b111010000100001100101111,
24'b111011000001111100000100,
24'b000011100111110111011001,
24'b111011100010000011001101,
24'b001011010010000101011110,
24'b111100100000110110110000,
24'b111010110111001110100110,
24'b111100001100111000011001,
24'b000111001001110110011110,
24'b000111010111000110011000,
24'b101111110010001000010100,
24'b001001011001111101000011,
24'b000000100000111001101001,
24'b111100110111111111000001,
24'b111101111010000010011011,
24'b000100101100001000011011,
24'b000000011000110111101101,
24'b111111011000000010101000,
24'b111010110000111001000001,
24'b000100110011000110110011,
24'b111101000011000100000010,
24'b000100111010111001111101,
24'b000001100100111111001111,
24'b110011001101111110010001,
24'b001100010111001010000101,
24'b111100000100110110010101,
24'b111011111010000011101010,
24'b000111010011111110000101,
24'b000100100010000011101110,
24'b101101101011111100101100,
24'b000111001111111101101110,
24'b001010111011001001101000,
24'b111010111000110111111011,
24'b111001100101111011111001,
24'b000001001110001010001110,
24'b000110000111111101101010,
24'b111010010000111011000111,
24'b000011011011000100111100,
24'b000000011010111001110110,
24'b111111010111000100101010,
24'b111011011000000010101000,
24'b000100000001111110111111,
24'b000000011000111000011100,
24'b000001010100000011100000,
24'b111110000110000101110111,
24'b000000000000111011000011,
24'b111110001011000101001001,
24'b111100101000110110011010,
24'b001100100010000100001000,
24'b111011101000000001011011,
24'b111001111000000111000101,
24'b111011111010110000111010,
24'b001011101110001100100111,
24'b111101011110111010110001,
24'b000000100101111000100101,
24'b111000110110001110011101,
24'b000111010101111110001011,
24'b111000011110110111000000,
24'b000100011100000000100010,
24'b001000000111000100010001,
24'b111000010001000001100100,
24'b111010110110000010100110,
24'b000010011101110111011101,
24'b000010100000000000100010,
24'b000110011101000101110010,
24'b000000100000111011110110,
24'b101111101000001000110010,
24'b111111110110110010001011,
24'b010011001100000111011001,
24'b111110100110000001100000,
24'b110111110011111011100010,
24'b110100010100000011001000,
24'b001001110001000000010001,
24'b001011100010000000000001,
24'b111001011111111101010010,
24'b111011110101111101011100,
24'b111100001011001010011010,
24'b111101010111110111101101,
24'b010011001100000011010100,
24'b111001100010111100001111,
24'b110111101111000011000100,
24'b110111101110000001100100,
24'b001101100000111010011001,
24'b001100011010000110100001,
24'b101011001010111100010111,
24'b000100100110000010100001,
24'b111101101010111010000100,
24'b000110000000000100101100,
24'b000110000110111110011101,
24'b110101110010000111101001,
24'b111100100011111000111101,
24'b000111001101110110000100,
24'b000001101011001011100100,
24'b111001111000001001110000,
24'b001001100110110001101000,
24'b110110110000111110010110,
24'b111000001100000010010101,
24'b010110100101001100000010,
24'b110100111111110010000101,
24'b110111110100000001001101,
24'b001010011110000111110001,
24'b111101110000000000100110,
24'b111010000011110000011101,
24'b001011010101001001111010,
24'b110111110100001000011100,
24'b000000111000111010100110,
24'b111110111011111000011001,
24'b000011011111000010010000,
24'b000010111101000010111100,
24'b110011100010000011110100,
24'b001111100110000001011111,
24'b110011111010110111001110,
24'b000100000111111010110110,
24'b000001101100001101000111,
24'b000100011001111111101111,
24'b101111001100111101111111,
24'b010000101001111010111000,
24'b111110010101111101000011,
24'b111000111101001001110111,
24'b111110111001111011010110,
24'b001000011110001000000010,
24'b111101111001110100011111,
24'b111110110000111101101010,
24'b110110100101001010110101,
24'b001100111010111100101100,
24'b000001100000000000000001,
24'b110111010100000001101100,
24'b111101001010111000101101,
24'b001001010111111111110011,
24'b111101111000001001001000,
24'b111111100010000011010010,
24'b111100010010110100101111,
24'b000011001001111110011100,
24'b111011011100000010100110,
24'b001011010001001000110100,
24'b111011101110111111100000,
24'b110001011011110101011111,
24'b001111011011111101010111,
24'b000001010101001101110010,
24'b111010111101111010110101,
24'b111011111010111111101111,
24'b000011001011111011011101,
24'b000100010001001000100010,
24'b111011100100110100110110,
24'b000010000010001001011100,
24'b111110111100111011000111,
24'b111111110100001011000101,
24'b111101000110101100101001,
24'b000101010001001011110110,
24'b000100010010111101000001,
24'b110010111010000100100100,
24'b000101110001111110000100,
24'b000011010110111101010010,
24'b111110011000111111001111,
24'b111110011010111111111001,
24'b000100100010000100010001,
24'b110111011011000001011101,
24'b000000111101111110101100,
24'b001101000101111000010110,
24'b110110011011111101001111,
24'b111111000001010101010111,
24'b111000011010101111011011,
24'b010010000101000110111111,
24'b110111100111111000011110,
24'b000011100011111010111110,
24'b101110111110010011010001,
24'b001111001001111000110010,
24'b000110111111111001011111,
24'b110110001001000001001010,
24'b111010010001000001000101,
24'b000101001010000010111110,
24'b000001100001111101101111,
24'b001001001010000111100111,
24'b110000111010110010111100,
24'b000011110010000010001000,
24'b111100110011000110110101,
24'b001101100101111110010111,
24'b110111000011111111110000,
24'b000000011000000000110111,
24'b111011000010111001100011,
24'b000100101100111111011101,
24'b000100110101001100010101,
24'b111100001111111100001011,
24'b111101001001111000100001,
24'b000001110101111111101110,
24'b111101110001001001011111,
24'b000100001000111000010100,
24'b000011101010000010010010,
24'b110100000100000011001110,
24'b001010000111111111110100,
24'b111010010101110100110110,
24'b000010000000001001100001,
24'b000010101111000001101110,
24'b111100010111000000110001,
24'b000000010011111010001010,
24'b000010110010111111001101,
24'b111011100101000001100001,
24'b000001001110000100000010,
24'b000100011100000010010111,
24'b111101010101110110010000,
24'b111110101110000100100111,
24'b111101000111000001101110,
24'b000101001000111011110101,
24'b000001001010000011110111,
24'b111011100011000010001111,
24'b000000111010111110000111,
24'b000101010000110110011110,
24'b110100010000001001110110,
24'b001000011110000001000111,
24'b000100111000111111010011,
24'b110111000010111100101000,
24'b000001110110111110001010,
24'b000010001000000000110110,
24'b111100010010000101110100,
24'b000010010111000001000111,
24'b000100000111110100111111,
24'b000001101010000110000001,
24'b110000110011000001111101,
24'b000101011110111111000010,
24'b001100000110111110000111,
24'b111010100000000000001101,
24'b000001101110000110000010,
24'b101110000011110011110101,
24'b010001110111001010011000,
24'b111110001111111101100101,
24'b000010011101111101001110,
24'b111000101100000011000000,
24'b000011110001111111111111,
24'b110111000101111101110001,
24'b001001010111111101101101,
24'b000110011000001000110010,
24'b111010011101111001001011,
24'b110110001000111111000011,
24'b000100100011000111000000,
24'b000100001100110111110111,
24'b000011010000000001010010,
24'b000010001101000111100010,
24'b110001111110111000101010,
24'b111101101010000101101001,
24'b010010000010110011111101,
24'b111110010111001101111110,
24'b110110000011111101110001,
24'b111101101011110100111000,
24'b000101101100010000001000,
24'b000101101001110100111010,
24'b110110001111111101001110,
24'b000110000111001100111000,
24'b000000101100110111110101,
24'b110011101011111110110110,
24'b010000110000000010010001,
24'b111011000010000000111100,
24'b111001010001000000001111,
24'b000010010011111100110111,
24'b000111100110111101001101,
24'b111010110011001101100010,
24'b111101101000110111011110,
24'b111110000001111000001000,
24'b001000101100000111100101,
24'b111110010101000001110110,
24'b111010000011000101110010,
24'b000010110111110100001110,
24'b111100011011111101100011,
24'b001001111100000111001001,
24'b111000101011000100101101,
24'b000001101100000000011110,
24'b111100101011110001001101,
24'b000011001110000110101001,
24'b000011110111000111000000,
24'b110011001101111101100000,
24'b010011101101111011111000,
24'b101111111001000010001111,
24'b000100100011111101100101,
24'b111001000010000101101001,
24'b010011011000111000010101,
24'b110011111010001000010100,
24'b111000111100111011000000,
24'b000110000111000000000101,
24'b000111110100000001011110,
24'b110110111111000000100011,
24'b000000111110110101100010,
24'b000010111010010110101101,
24'b111100011101110001011000,
24'b000100010000111000111110,
24'b111101011110000111011100,
24'b111011101110000110001110,
24'b001011101000111111110000,
24'b110101010110110001101111,
24'b000100100011001001011111,
24'b111011111111000011011101,
24'b000100110010111011011101,
24'b000000001010111100010100,
24'b111111100011001011110110,
24'b111001010011110100010010,
24'b000100110011000011001110,
24'b000111110001000000111111,
24'b110100010000000001100011,
24'b000010111110000000101000,
24'b000010000100111001001111,
24'b000011011111000111110001,
24'b111001110010111101111000,
24'b111111000111110111011011,
24'b000010111101001110011000,
24'b000101110100111010111101,
24'b111100100000111101111011,
24'b110001100010111001011100,
24'b010010100000000101100001,
24'b111101001010001010000001,
24'b111011000011111110110110,
24'b000010100010100101101010,
24'b111001001011010110010001,
24'b001000000010000011110110,
24'b000100110010111011111111,
24'b110010011000110101100100,
24'b001000110010000101100000,
24'b111100100000000100001110,
24'b000000010111111110111110,
24'b000111001001000001010100,
24'b110101010011111000001110,
24'b000010111010000000011011,
24'b000011110111001111100101,
24'b000000101101110001110010,
24'b111001111111111101111011,
24'b000001110101000110010100,
24'b000001110110000010101100,
24'b000100000110000000010111,
24'b110111100101110010111101,
24'b000011100001000110101111,
24'b000000101000001011111011,
24'b111100110101110011111000,
24'b001100110010000011010000,
24'b101110110100110111110100,
24'b000010001101001000001110,
24'b001100001101001001100101,
24'b111011100111110000010010,
24'b111000010001000000001111,
24'b000010100011001010010110,
24'b000110001101111000010011,
24'b111110011010000000101011,
24'b111010101010001001101011,
24'b000010110100110011011000,
24'b000000011110000010010010,
24'b000001111010000000110000,
24'b111100001001000111101001,
24'b000100110010111000100110,
24'b111000110011000101111100,
24'b000101011100110000110110,
24'b111111101000001100110110,
24'b000010000100000010001111,
24'b111010110000000000000110,
24'b111110011101110101101101,
24'b000111110101000010010001,
24'b111110111000000100110001,
24'b111000101001000011000010,
24'b000111101011111110110111,
24'b111001100100110100100110,
24'b000101011001001110100010,
24'b111111111110110000110000,
24'b111010001011010001001111,
24'b000111011100111010001110,
24'b111001011111111001111111,
24'b000101100011111101101010,
24'b111001101100001100100011,
24'b000110010001111001011101,
24'b000001001101111110100011,
24'b110101000010000001011010,
24'b001001110010000000100101,
24'b111111001000111110100001,
24'b111110010101000000101100,
24'b111101010010111110101100,
24'b000110100011000111110100,
24'b110111111111110111101110,
24'b000110010000111011011110,
24'b111111010000001000100001,
24'b111101111011000011110111,
24'b111110010010111100010010,
24'b000011010100110101000111,
24'b000100010101000100000111,
24'b110110111100010011100011,
24'b111110111111110001000100,
24'b001010101101110000001000,
24'b111011110010010111001100,
24'b111110111110000010000111,
24'b111000011010101101001101,
24'b001001000001001000101111,
24'b000000111000000110100110,
24'b000001111101110101000011,
24'b110101010010000100011000,
24'b000011001101001000111001,
24'b000011000010110001000001,
24'b000110101010000100111101,
24'b110111001000000100011101,
24'b000000010000000000101100,
24'b111111111100111000110011,
24'b111111000111000100101000,
24'b001000001000000001101100,
24'b111111010100110110111000,
24'b110110000010001100101110,
24'b111100111101111000111101,
24'b001111100010000010100000,
24'b111100001111111101101110,
24'b111100000000111000010001,
24'b111100011101010001011011,
24'b000010111000111010011101,
24'b000001001010110111010111,
24'b000100110111000011101010,
24'b1_11100100101111111010111,
24'b111110001010111110111001, 
24'b000100111110111011110111, 
24'b110111000110000110101100, 
24'b000100101111111100000111, 
24'b000101010010111110111011, 
24'b110110101001000011110100, 
24'b000011100011111100110110, 
24'b000011101101000000101011, 
24'b111010110101000001011010, 
24'b000001110011111110011101, 
24'b000011110111000000010110, 
24'b110110011100111111101110, 
24'b001000010010000010010010, 
24'b000101010000111100100101, 
24'b101011100101000001000010, 
24'b010010101010000010110010, 
24'b111111001011111011101010, 
24'b110110010111000100011110, 
24'b000000101000111001100101, 
24'b001000111011001000001100, 
24'b000010000111111100001101, 
24'b101001001111111010000001, 
24'b011001100101001011011010, 
24'b111000000001111000111111, 
24'b111010100101000000011101, 
24'b000001010010111110100000, 
24'b000110001100000111001000, 
24'b111101110011111001101010, 
24'b111010000111111101100011, 
24'b000100100110001000011100, 
24'b000011100110111011101101, 
24'b111000010010111100011111, 
24'b000111100001000101010001, 
24'b110101110001111110101001, 
24'b001110111011111111001011, 
24'b110010010001111110101011, 
24'b000110100011000100001111, 
24'b111101011000111010000111, 
24'b000110100110000111100111, 
24'b110010111011110111110001, 
24'b001111010000000011110111, 
24'b110011110001000100011110, 
24'b000110101011110110011100, 
24'b111110110010001000000110, 
24'b111110100010111001100001, 
24'b000000101000001011100110, 
24'b000000011101101101000101, 
24'b000001110110010001010100, 
24'b111010001101111010101110, 
24'b000110101001111010111001, 
24'b111100010000000011100111, 
24'b000000000001000100100110, 
24'b000011110001111001101110, 
24'b111000000000111110101110, 
24'b001001000010000111000111, 
24'b111101001011111101100000, 
24'b111010000001111001100001, 
24'b000111100100001000001000, 
24'b111110110011111110001010, 
24'b111101001010111111001000, 
24'b111111100011111001001000, 
24'b000010011100010001000001, 
24'b000100101111101111000110, 
24'b110010011101000101110001, 
24'b001011011101000100011001, 
24'b111111011101111100000111, 
24'b111011001000111011100111, 
24'b111111100001001010000010, 
24'b000110001101111000100101, 
24'b111101000001000000001001, 
24'b111100100011000100111011, 
24'b000010010110111011000101, 
24'b000101000111000010101110, 
24'b111000101100111101110001, 
24'b111111110011000011010010, 
24'b000111010011111110000011, 
24'b111101100101111100011100, 
24'b110100101101001001001101, 
24'b010010101111110101101101, 
24'b110100101001001001000111, 
24'b111101101000110011111101, 
24'b000111111111010011000001, 
24'b111100111001101011001011, 
24'b111110100010001011011010, 
24'b111110000011000010010011, 
24'b000111110011110111100111, 
24'b111001100010000100101100, 
24'b111110010101000001001110, 
24'b000111011101111011001110, 
24'b111010100010000111111101, 
24'b111111000101110110011101, 
24'b000110000011000011000101, 
24'b111000010011001010100001, 
24'b000110100000101110011010, 
24'b111011011101001000100011, 
24'b000101100001000110000011, 
24'b110101000110110111111110, 
24'b001111110110111101000010, 
24'b110010100110001001101001, 
24'b000011111101111100001001, 
24'b000100100010111110010101, 
24'b111000110110111011001110, 
24'b000111010100001110000010, 
24'b110111010111110110001010, 
24'b000111110110111011010101, 
24'b111110111011001011000010, 
24'b111000110000111100101011, 
24'b001001000111111011100101, 
24'b111011111001000001100100, 
24'b000000001111000011010101, 
24'b111101010111000000110110, 
24'b000111100110111000000011, 
24'b111000001010000100110101, 
24'b000001011101000110000101, 
24'b000110100010110110101001, 
24'b110111000001000000111110, 
24'b000011100100000110001111, 
24'b000100001001111100010000, 
24'b111010101100000000001101, 
24'b111101111110111011001111, 
24'b001001101010001010010110, 
24'b110111001011111010010111, 
24'b000000111000111011110100, 
24'b000101100011000011111111, 
24'b111001111011000110101100, 
24'b000011111001110100011111, 
24'b111101110110000010111110, 
24'b000000001101000101110000, 
24'b000001111111111101101011, 
24'b111110011100111011011101, 
24'b111110010000111111110011, 
24'b000011001110001011101100, 
24'b000000010000110101110000, 
24'b111011010101111000001100, 
24'b000011110000010110001011, 
24'b000010101000110000011100, 
24'b110111110111111100001101, 
24'b000110110001001111110110, 
24'b000010000110110001111010, 
24'b110011011000000110111000, 
24'b010000001111111111011110, 
24'b110110110110111010101110, 
24'b111101111101001000001001, 
24'b000110001010111101011101, 
24'b111111111111110111100010, 
24'b110111100100001100110001, 
24'b001011011011111010111011, 
24'b110110111000111011010001, 
24'b000100001101000101010100, 
24'b000011101010000001111100, 
24'b110011111110110111110001, 
24'b001100100110001011000101, 
24'b111101100100110010000011, 
24'b111000001010010000100001, 
24'b000111110111110001101101, 
24'b111100011111000111110001, 
24'b000110101000111100111000, 
24'b110011100010000011100001, 
24'b000101100011111001111010, 
24'b001100001100001000100010, 
24'b101101000110110100110110, 
24'b000101100011001011011011, 
24'b001000001100111011100101, 
24'b111100000111111000100011, 
24'b111001011101001100011111, 
24'b000001000111111100000001, 
24'b001111010011110110010001, 
24'b101110000100001111100011, 
24'b000010111100110100000100, 
24'b000101011010000111011110, 
24'b000110101011111001100010, 
24'b101011100001000100110010, 
24'b001110000000000000001101, 
24'b000101010000111011011011, 
24'b110010000111000101000010, 
24'b000110111111111100010010, 
24'b000000010110000010101111, 
24'b111111110111000000011001, 
24'b111111111111111000111000, 
24'b111011111100001100100101, 
24'b000100000111110100111111, 
24'b000100000100000011100011, 
24'b110110000100000011110100, 
24'b000011111010111000100011, 
24'b000101111111000111010101, 
24'b111010111111111011101011, 
24'b111001101110000000100010, 
24'b001101100001111111011101, 
24'b110101110111000110100110, 
24'b000101110001110010010110, 
24'b110101110000001110101100, 
24'b010010011001110101110111, 
24'b101110100100000110000011, 
24'b000100101001111011111101, 
24'b001001100001000000100110, 
24'b110001111000000010110001, 
24'b000111110011000001101010, 
24'b000010111001110010101101, 
24'b110110000100010001100000, 
24'b000111101101111100011010, 
24'b000011101011101111011000, 
24'b101111101101010100011001, 
24'b010011101010111100000100, 
24'b110100000000110100010111, 
24'b000011101011001000001100, 
24'b111011100101000110110001, 
24'b001010000000110010101101, 
24'b111000001100000110111010, 
24'b111010111000111111000010, 
24'b010001001011000100100110, 
24'b101110101101110101100111, 
24'b001000001100000111111010, 
24'b111111111010000000100101, 
24'b111100011001111010111110, 
24'b000110101111000010111011, 
24'b110110000011111111011110, 
24'b001000110111000001010100, 
24'b111101000100111111001010, 
24'b111111001010111011100000, 
24'b111101011011001010010101, 
24'b001000101110110110010110, 
24'b110110111000000010101111, 
24'b000010101000000011010101, 
24'b000011010111111100010000, 
24'b111101111010000000111111, 
24'b111010111011000000011000, 
24'b001011000101111111011110, 
24'b110100111011000011011101, 
24'b000110111111110101111011, 
24'b111100010111001111011101, 
24'b000010011001110010000011, 
24'b111111100100000110010010, 
24'b111100111001000001001010, 
24'b000100000111111100100011, 
24'b000000010110000010001100, 
24'b111010001001111110000001, 
24'b000110000010000100011111, 
24'b111110001111111000010100, 
24'b111111001110001001100111, 
24'b000000110110110110010011, 
24'b111100010111000111000111, 
24'b001000111010111110010101, 
24'b110111011000111100110101, 
24'b000000010010000010110110, 
24'b000110001101000001010101, 
24'b111101101011111101110000, 
24'b111010011001111100101110, 
24'b000110011111001000111100, 
24'b111101110011111000100110, 
24'b000011000100000001011110, 
24'b110111000010111111111001, 
24'b001000101100000101011011, 
24'b000000110100110101011011, 
24'b110111110100001010100001, 
24'b000101010001111000101100, 
24'b000001000111000011111100, 
24'b111110001010000000011000, 
24'b111111101000111011010101, 
24'b111110101110000100100000, 
24'b000100100110111111111111, 
24'b111100010000111111000111, 
24'b000001101101111010101111, 
24'b111010101011001001010100, 
24'b001011010001111101111001, 
24'b110110101101110111000110, 
24'b111111100000001000110101, 
24'b000101110011000001000001, 
24'b000000010010111101000101, 
24'b110110100011110101110110, 
24'b001011000001010101110110, 
24'b111010100011110000110011, 
24'b000000101110111101100101, 
24'b111110110001001001101100, 
24'b000101110001111111011101, 
24'b110101010001110101011100, 
24'b001011011110001011010000, 
24'b111011010101111010100010, 
24'b111010011111000010101110, 
24'b001001000111111100011001, 
24'b111101010001000010111000, 
24'b111100000000000000001111, 
24'b000001001010111110100011, 
24'b000111001011111110100010, 
24'b110111001110000101111010, 
24'b000001000100111000000011, 
24'b000101011101000101110110, 
24'b111101111001111110101000, 
24'b111001001000111111001000, 
24'b001011001101111101100101, 
24'b111000110011001000000010, 
24'b000000110100110111100111, 
24'b111111110000000000100110, 
24'b000111000111001001010011, 
24'b110001101101110010101001, 
24'b001101011010001010001001, 
24'b111011001000111100010110, 
24'b111110010010111101110011, 
24'b000000011100000100110111, 
24'b000010111110111110000110, 
24'b111111001011111010101001, 
24'b111100111000001010101011, 
24'b111111001110110110101001, 
24'b001010110101000100110100, 
24'b110010011101111101001010, 
24'b000010111001000010000010, 
24'b001010011011000011001000, 
24'b110010001100110101110110, 
24'b001000001010001001101101, 
24'b111110000001111111001110, 
24'b111110111000111011110100, 
24'b000001101011111100010010, 
24'b000001110110001111011110, 
24'b110111011101110001001001, 
24'b001010100001000000101001, 
24'b111101001000001011111100, 
24'b111010101100110100010111, 
24'b000010011100000011111101, 
24'b000110011110111111010010, 
24'b111001111001000011100110, 
24'b111011111101111011100000, 
24'b000111001011111110101110, 
24'b000100000100001000011110, 
24'b110001111000110111101110, 
24'b000111110011111110101100, 
24'b000101111010001101101100, 
24'b111000010010101100010000, 
24'b111101010001001111100011, 
24'b001000000000111011001100, 
24'b000000010101111011011010, 
24'b110100101000000110111111, 
24'b001101101100111101010101, 
24'b110101111011111101010010, 
24'b001000110111000010111011, 
24'b110101010111000011100100, 
24'b001010101000110100011010, 
24'b111000101011001101000101, 
24'b000010110101111010111111, 
24'b000001000101111001000100, 
24'b111110000011001101111001, 
24'b111101010111110011000101, 
24'b001001010100001001010011, 
24'b110111000101110111001000, 
24'b111110111001001011001101, 
24'b001010101001110100111111, 
24'b110110001101000101111101, 
24'b000010111001000000000001, 
24'b111111011011111110100101, 
24'b000010001010111110001101, 
24'b000001111101000011000101, 
24'b110100111011000011001110, 
24'b001011110110110010001001, 
24'b000000100101010010001000, 
24'b110100000100110110001111, 
24'b001000110111111100010011, 
24'b000001000100000111101101, 
24'b111110000001000010101000, 
24'b111011011011110000001001, 
24'b000010101000010001011110, 
24'b001010111110111001001111, 
24'b101101001110111100011010, 
24'b001000100101000011101101, 
24'b000111101110000010101000, 
24'b110100111100111010111011, 
24'b000001001111000000010000, 
24'b000110110001000101111100, 
24'b111001011011111000100010, 
24'b000101011011000101001010, 
24'b111000110010111100110010, 
24'b000110001101000010111001, 
24'b111111001011111101011110, 
24'b111111111001000010000110, 
24'b111000110101111100000011, 
24'b001011011011000111111101, 
24'b111101001010110110100110, 
24'b110110101001000100101110, 
24'b001000100011000011001101, 
24'b000100110001111000000001, 
24'b110001110101000111100011, 
24'b001011101001111010110000, 
24'b111001110111000100001100, 
24'b000101111001111011111100, 
24'b111001001110000011110111, 
24'b000100011000111100010011, 
24'b111011111110000010101110, 
24'b001001100000000000110100, 
24'b110100000110111011000101, 
24'b000010011111000100000110, 
24'b001010110111000011010000, 
24'b110011001111110100111000, 
24'b000010101001001110001100, 
24'b000101110110110001001111, 
24'b111010011010010000001000, 
24'b000010101100110010101101, 
24'b111101101010000000000011, 
24'b000001010010010000110001, 
24'b000001101011101010011010, 
24'b111111000111001010101011, 
24'b111011011110000010000100, 
24'b000101100000111011100000, 
24'b000010011111000001110000, 
24'b110110100010111100000001, 
24'b000101010111001000011110, 
24'b000100010000111010101100, 
24'b111001001011111100101111, 
24'b000001010101000100000000, 
24'b000011101110000110101011, 
24'b111010010011110000100010, 
24'b001000001010001010010110, 
24'b110110111000000011110001, 
24'b000010011101110011000010, 
24'b001000100110001011011000, 
24'b110010110110111100000011, 
24'b001001011011111101110011, 
24'b111000101001000010101011, 
24'b001010011110000011110111, 
24'b110111001000110010111011, 
24'b111100111001001111101010, 
24'b001111000010111000111100, 
24'b110000110000111011011011, 
24'b001000000011000110111011, 
24'b111011011010000000110101, 
24'b000100111000111000111000, 
24'b111111010010000011110001, 
24'b111000011001000100001001, 
24'b001011000001111001100101, 
24'b111001111110000000111000, 
24'b111110100010000110001101, 
24'b000110101011110111001001, 
24'b110110000000000110100011, 
24'b001010110001111101100111, 
24'b111001110111111111111010, 
24'b111110011101111110111111, 
24'b000101010111000100011111, 
24'b111100100101111010000001, 
24'b000000100000000010010011, 
24'b111111111111000100011000, 
24'b000001000010110111001100, 
24'b111101001010001000101111, 
24'b000100001100111000111001, 
24'b000000010101000111010100, 
24'b110100000110110111010010, 
24'b010001010110001000001010, 
24'b111100111011111010111011, 
24'b101100101101000010000111, 
24'b010101000000111110111011, 
24'b000011011101000000100110, 
24'b101000011010000000110110, 
24'b001110100010111110001010, 
24'b000111101001000000100011, 
24'b110100010001000001001011, 
24'b111101110110111111110100, 
24'b001000111000111101011101, 
24'b111110010011000010101011, 
24'b111111010100111111111010, 
24'b110111011010000000011100, 
24'b001011011011111001111110, 
24'b000001111100001010001010, 
24'b110011011010111010000000, 
24'b000010000000111101010100, 
24'b010011000011000101111010, 
24'b100011111011111110011101, 
24'b010110100001111100111001, 
24'b110001100010000011010010, 
24'b000110101110111101011000, 
24'b000101100000000100000010, 
24'b101111100010111100010010, 
24'b001110111110111110111110, 
24'b111100000100000100111110, 
24'b111100101000111101100011, 
24'b000100001101111101100000, 
24'b111001111110000010000011, 
24'b000111101110000011100000, 
24'b111111001110111001000010, 
24'b110101010111000110000011, 
24'b001011001101111010101011, 
24'b000000000111000110100110, 
24'b111010010111111010110000, 
24'b111101010010111111011000, 
24'b001010000110000101001110, 
24'b111100111001111100111011, 
24'b110110100000111110000100, 
24'b001101011010000001001101, 
24'b110110000000000111110110, 
24'b000111011110101110000001, 
24'b111011100111010011001000, 
24'b111101110011110111100101, 
24'b000100100011111010100110, 
24'b000010001101001000111011, 
24'b111010111110000000100101, 
24'b110111010101110110011111, 
24'b011001100011000011111100, 
24'b101001101010001010011110, 
24'b000010000000110010000000, 
24'b001001110111000000101111, 
24'b111100010011001011011110, 
24'b111100000011111010100011, 
24'b000010000100110100111001, 
24'b111111100110010001010001, 
24'b000101001011111000001010, 
24'b111011110100111100111110, 
24'b110111010111000100101001, 
24'b010000000110111110011001, 
24'b111011110111000001010111, 
24'b110100011101111101010101, 
24'b000111100001000010001010, 
24'b001010101001111101111101, 
24'b101110111000000100100011, 
24'b000100001111111010101110, 
24'b001010100101111111101101, 
24'b110010010000001000110111, 
24'b001001110110110010100010, 
24'b111010011100001100011001, 
24'b111111101000110111100010, 
24'b000110111100000011010010, 
24'b111000110101000010010110, 
24'b000000011100111010011010, 
24'b000101000100000100110101, 
24'b111010000011111011111100, 
24'b000111010001000111101001, 
24'b110111000100110011110011, 
24'b000100000010001001110000, 
24'b000101010111000001000111, 
24'b111001100000110100001100, 
24'b111101010100001101010000, 
24'b000111101001111010110000, 
24'b111110101100111011110011, 
24'b111101011010000111011011, 
24'b111001101000111011100000, 
24'b001111101001000010000000, 
24'b110101110011111100000110, 
24'b111111100100000100110100, 
24'b111101111101000010101001, 
24'b001101000000110001110100, 
24'b110011101011010000001111, 
24'b111110111111111010100010, 
24'b000110111011111100000111, 
24'b000010101110000000011101, 
24'b110011101000000110010010, 
24'b001001011101111111000001, 
24'b111110110110110100100010, 
24'b111100111000001100110001, 
24'b000110011000111110101100, 
24'b110101011000111011111101, 
24'b000111001110111010110110, 
24'b000110001101001100101100, 
24'b110001111000111011001110, 
24'b000100011100111001010101, 
24'b001010101110000100001001, 
24'b110100000011000101111001, 
24'b000001011010111100101001, 
24'b000011100111110100101100, 
24'b000001001110001111110000, 
24'b111100001001000000110001, 
24'b111110110010101010111111, 
24'b000101111100010111100010, 
24'b111011000111110111011111, 
24'b000011000010111001000101, 
24'b111100100101001010000011, 
24'b000001110000111110100010, 
24'b000011010001110110010011, 
24'b111010110101001101011110, 
24'b000001000111111001110100, 
24'b000011010001111011010001, 
24'b111011111010000111101100, 
24'b000100110010111111000100, 
24'b111001000101111001111110, 
24'b000110010011000110110100, 
24'b111101000101111010100110, 
24'b000011101101000110010010, 
24'b110110001100111001100001, 
24'b001100001001000011110100, 
24'b111001011011111100110011, 
24'b000010100010000111011110, 
24'b111001010101110110010100, 
24'b001001101111000100010101, 
24'b111110101011000001010101, 
24'b110100110110000010001001, 
24'b001101000001110110010000, 
24'b111011010001001001000010, 
24'b111110110011111111110110, 
24'b000001101010111011001111, 
24'b111011101010000001100000, 
24'b001010001111000001000001, 
24'b110100100010000010110110, 
24'b000111100111111001100111, 
24'b111000111001000011001010, 
24'b001001110110000010110101, 
24'b111011100010111011001001, 
24'b110101010111000010111100, 
24'b010100010110000000011010, 
24'b110000110110111010000100, 
24'b000101100110001100100001, 
24'b111101000010110001110001, 
24'b000000100000001000110010, 
24'b001010100001111101100001, 
24'b101101010100000000010101, 
24'b000111011000000010000000, 
24'b001111100011110110111111, 
24'b100111011000001111110000, 
24'b001101011010110000010111, 
24'b111101010101001011110110, 
24'b000111010000110100100011, 
24'b110000101010001100100100, 
24'b001011010111110111010100, 
24'b111101111100000001111111, 
24'b000011110001111111111010, 
24'b110001101010000001111101, 
24'b010000101010000000111011, 
24'b111010001010110111011101, 
24'b111011110001001010110101, 
24'b000011110111111011101110, 
24'b111110101000111110001111, 
24'b000111010111111111110100, 
24'b101111011100000101011011, 
24'b001111001000111000101100, 
24'b111111001100000111001010, 
24'b110001110111111001000101, 
24'b010010101011000010001101, 
24'b110001110101001001000101, 
24'b001000011110101101110100, 
24'b111010101111010000101000, 
24'b000010111100110110100011, 
24'b111111101011000111100111, 
24'b111111000111110101001110, 
24'b111110111110001001011000, 
24'b000101100011111110111111, 
24'b110101100001111001111110, 
24'b001101001101000110000011, 
24'b110101000101111101000010, 
24'b000011010100000010001001, 
24'b000101010111111100001100, 
24'b110111101010000110100110, 
24'b000011010000110110100010, 
24'b000101101010001000111110, 
24'b110011111010111110010110, 
24'b001101010001111000011101, 
24'b110110110101001000011110, 
24'b000000100101000000001001, 
24'b001001000010111001010101, 
24'b110011011100000010011111, 
24'b000110000111000110000000, 
24'b000100001111111000010111, 
24'b110111111011000010110001, 
24'b000011011101111111010001, 
24'b000001011110000100111001, 
24'b111111110100110111100111, 
24'b111011000100000100110100, 
24'b001000100101000011101011, 
24'b110110010001110101110100, 
24'b001000101110001010101100, 
24'b111100010000111001010010, 
24'b111011110011000011011011, 
24'b001000001000111010111000, 
24'b111100101000001001110111, 
24'b111100000001110101101000, 
24'b000101000101000011001110, 
24'b111111000001000100110101, 
24'b111111101010111011100000, 
24'b111101101101111100100101, 
24'b000010100000001000110111, 
24'b000000100000111010001111, 
24'b000001001010111111101011, 
24'b110101101101000000110010, 
24'b010001011001000100100110, 
24'b110010011111110111110100, 
24'b000011110000000100001111, 
24'b000001000111000011111010, 
24'b111111101110111000111110, 
24'b000010010101000000001100, 
24'b110101111010001010111010, 
24'b001111110110110001010100, 
24'b110011111011000111000100, 
24'b000001100100000011101011, 
24'b000110011000111000100101, 
24'b111010010100000100100010, 
24'b111110011010111101101010, 
24'b000111111010000011001011, 
24'b111001001110111100111111, 
24'b111111010101000001100111, 
24'b000101101100111011111110, 
24'b111111010101001010011100, 
24'b110100010000110010111011, 
24'b010100011110000111101110, 
24'b101110101111111111100000, 
24'b000100011000111101101110, 
24'b001000101100000011111111, 
24'b110010001100110110010100, 
24'b001010011100001110110111, 
24'b111011010100110100100010, 
24'b000010110001000001100100, 
24'b111011011000000101001110, 
24'b000101111001111010010010, 
24'b111010011100000101011010, 
24'b000111000111111001111010, 
24'b110110000100000010101000, 
24'b000110111111000110000000, 
24'b000011101001110101000101, 
24'b110100110110000101001011, 
24'b000110000010000101101001, 
24'b000011100111110110111000, 
24'b111101101000111111100110, 
24'b111000100110010001101111, 
24'b000111001110100000110110, 
24'b001000000010011110010100, 
24'b101100111111110001011011, 
24'b001010000000111101001110, 
24'b000110011110000101110000, 
24'b111000000001000101000101, 
24'b111011011110110100101100, 
24'b001010011001000000110101, 
24'b111110000111001111000111, 
24'b111010101001101110011101, 
24'b111101110001000110001001, 
24'b010000010010000010101011, 
24'b101100010001111111001111, 
24'b001001001110111101011011, 
24'b000100000100111110010110, 
24'b110110010011001000101110, 
24'b000111001101110101110011, 
24'b111100110110000110110101, 
24'b000011101101111100110010, 
24'b110111110111111110010101, 
24'b001000110111001001101101, 
24'b111110001101110000111000, 
24'b111011010010001011000101, 
24'b111111001011111110011000, 
24'b001110110001111101110011, 
24'b101100000011111101110111, 
24'b001001100110000110011000, 
24'b000010100101111011010101, 
24'b111101010010000000101001, 
24'b111100100110000001001011, 
24'b000010000100111101111110, 
24'b000110010110000011100001, 
24'b110101000011111101100100, 
24'b001001110110111100110101, 
24'b110101001011000111111001, 
24'b001110101001111010010100, 
24'b110011100100111111001010, 
24'b000010000010000100010110, 
24'b000110101111111100100010, 
24'b111001010100000010111100, 
24'b000010000011111100010010, 
24'b000001100100000001011101, 
24'b111010110110000100011111, 
24'b001001110001110111110111, 
24'b110100011001000111000100, 
24'b001001010001111000011010, 
24'b111001010101001110110001, 
24'b000100101011101001111110, 
24'b000000110001010011000100, 
24'b111001010100111000111011, 
24'b000010011111111101100101, 
24'b001010111101000011111100, 
24'b110000111100111100010000, 
24'b111111111111000111001011, 
24'b010000010000110110110011, 
24'b110100000001000100010101, 
24'b111011110001000001100000, 
24'b000110011001000001100111, 
24'b000111001101110101001001, 
24'b110100100011001100111000, 
24'b111100100000111100101110, 
24'b001110111101111010000110, 
24'b111011111101000011000101, 
24'b110010011010000111000100, 
24'b001101000000110100101101, 
24'b000001100110000110011100, 
24'b111001110000111110111001, 
24'b111100000001000001001010, 
24'b001011000001111100100110, 
24'b111001111101000100010101, 
24'b000001001010111010001100, 
24'b111011100010001000011011, 
24'b000101010101111001100010, 
24'b000100101110111100111110, 
24'b110010101100001011110000, 
24'b000100100110110110100000, 
24'b001111001110000000100010, 
24'b100110011110000000001101, 
24'b010010110001001010111101, 
24'b111001101110101101111011, 
24'b111110011111000111001010, 
24'b000101111010001100001100, 
24'b110111011000101110001000, 
24'b000100100101000101101100, 
24'b000111011011000101010101, 
24'b101111110111111110111000, 
24'b001010100100111000000000, 
24'b000011010101000110011000, 
24'b110111011010000000101000, 
24'b111111110110000100010000, 
24'b001001110100101100101101, 
24'b111001100010010110101010, 
24'b111001111011111010000011, 
24'b001100000101110101100100, 
24'b111011011101000111000001, 
24'b111001000010000101111001, 
24'b001001111001111010010100, 
24'b111011111100111000111100, 
24'b111111110011001011111010, 
24'b111100100010111100110110, 
24'b001001101100111101100001, 
24'b110111010010111011100111, 
24'b111110110001001010100100, 
24'b001011011000111011011000, 
24'b110100010110111101000101, 
24'b000001110110111110111111, 
24'b000111110110001000000011, 
24'b111000011100111101010010, 
24'b111110101011110110110011, 
24'b001000011001001000000110, 
24'b111001011010000111010100, 
24'b111111110001101110111001, 
24'b000011111111001010011100, 
24'b111101100101000001000010, 
24'b111111101011111011101011, 
24'b000000101111000010011111, 
24'b000001010100111101100101, 
24'b111011001100000001100110, 
24'b000111111101000010101001, 
24'b111000111000111100000001, 
24'b000001010001111111100011, 
24'b000011010010000000101001, 
24'b000000100101001010001001, 
24'b110111011000101100100011, 
24'b001000111010001100011111, 
24'b000000011010000011010100, 
24'b111001011000110111110001, 
24'b000001011101000000111000, 
24'b000101010101000010000100, 
24'b111110111000000100101001, 
24'b110111000100111001010001, 
24'b001010001100111101100111, 
24'b111110001100000111001110, 
24'b111100101111000100101011, 
24'b000000111011101100000001, 
24'b111111110001010010100100, 
24'b000011001010111100001001, 
24'b000001111111111100010111, 
24'b101110100100111101101101, 
24'b011000001001000111100000, 
24'b110111100100111101001010, 
24'b110011001000111101101000, 
24'b001101000111111101101011, 
24'b000101110001001011011011, 
24'b101111110101110011010010, 
24'b000101010000000101010100, 
24'b001010010010000000101001, 
24'b110010111111000001010010, 
24'b001000000110111000101101, 
24'b111001001001001010010101, 
24'b000101111010111000001001, 
24'b000010011011000010110010, 
24'b110100100000000000110001, 
24'b001001011110111110110011, 
24'b000000000110000001100001, 
24'b111100000001111001110001, 
24'b000001010111001111011010, 
24'b111101000100101001101010, 
24'b001001010000010100000110, 
24'b110111011010110110100010, 
24'b111110111011111110111111, 
24'b000110001010000100010110, 
24'b111111100000111110001100, 
24'b111101101101111111110110, 
24'b110111101000111111000111, 
24'b010011110010000000110110, 
24'b110010001100000011011000, 
24'b111100010110111001000101, 
24'b001001111101000010011101, 
24'b000001111100000111110100, 
24'b110000000001110011011010, 
24'b010010101110000110010101, 
24'b110001001111000010110110, 
24'b001100100110111011001000, 
24'b110101001110000001111101, 
24'b000101111001111101000111, 
24'b111101110001000111101010, 
24'b000011001010110111100111, 
24'b111101011110000100001101, 
24'b111011111101111101010111, 
24'b001000100011000100111111, 
24'b111100101100111101010001, 
24'b111101010111111001111110, 
24'b111011010101001001010111, 
24'b010011011001000000010000, 
24'b101011011111110101001001, 
24'b000010111110000111001110, 
24'b001100110101000101001110, 
24'b110111010111111000011101, 
24'b110111111101111011100010, 
24'b010010001011001110100100, 
24'b101111001001110101101000, 
24'b001101000111111111100000, 
24'b110100101010000011110111, 
24'b000111011011000010111000, 
24'b000000000000110100011001, 
24'b111001011011001111001000, 
24'b001010010000110100101010, 
24'b110011100111000010011100, 
24'b001010111111000100110101, 
24'b111101001010111100010101, 
24'b111001000010111100010110, 
24'b001000001010000111001010, 
24'b111111111101111100111011, 
24'b111001011010111111100100, 
24'b000101101001111101000101, 
24'b111100011010000110111000, 
24'b000110111100111100000110, 
24'b110100111011111110100010, 
24'b001001010100000000110010, 
24'b111011100001000010111011, 
24'b000010111001111111001011, 
24'b111100001010111011010010, 
24'b000011110100000011010000, 
24'b111010101001000100101100, 
24'b001011000101111001111011, 
24'b110001110100111100100101, 
24'b000111001110001011001101, 
24'b000010111100111001101101, 
24'b111101001110111010110010, 
24'b111001011000001011100011, 
24'b001010101111110100010111, 
24'b111010001111001011100001, 
24'b000101010001110100011010, 
24'b101111110111001000011000, 
24'b010111101111111100010010, 
24'b110010111001000010101001, 
24'b111001101010111011100100, 
24'b001100111101000100111011, 
24'b111101010101111011000111, 
24'b110111011111000111111010, 
24'b001001100100110101000010, 
24'b111010011111000111000101, 
24'b000010111001000010110101, 
24'b000000110101110110011101, 
24'b111000011100001000101100, 
24'b001010101100111010001111, 
24'b111011011000000101101101, 
24'b111011000010111010111111, 
24'b001000101011111111001111, 
24'b111010010111000111100100, 
24'b000001011110111001110000, 
24'b000001011110111010001101, 
24'b111011110011010100011000, 
24'b000101010010100111010101, 
24'b111101100101001100100010, 
24'b111110100110001000001001, 
24'b000000101110101011100111, 
24'b000011001110001111000111, 
24'b111100101001111110011001, 
24'b111101100111111011110011, 
24'b000111010000000000101110, 
24'b111011000101111111111010, 
24'b111110010000000111000101, 
24'b000101011110110101000110, 
24'b111011101010000100001100, 
24'b000010011101000010110010, 
24'b111101000111000001111111, 
24'b000011110011110100110101, 
24'b111101101101001000000101, 
24'b111110110011000110101111, 
24'b000100010000110001010100, 
24'b111010100011000110100110, 
24'b000100111110000100010000, 
24'b111101000111111101111100, 
24'b111111011011110101111011, 
24'b000011011000010001000001, 
24'b111100101100110011100100, 
24'b000001111101000011110011, 
24'b111100001001000000011100, 
24'b001000111010111111110110, 
24'b110110010110000000011000, 
24'b000000110110111100101100, 
24'b001010110101000101010100, 
24'b110010011010111110111011, 
24'b000110011111111000000110, 
24'b111111001111001011011110, 
24'b000010111000111101110100, 
24'b111010010011110011111101, 
24'b000001011101001111000000, 
24'b000101001010111100011100, 
24'b111010101100111001000110, 
24'b000001011010000100000011, 
24'b111110000000000100011000, 
24'b000101101110111100011111, 
24'b111101010100111010000110, 
24'b111000010110001010110111, 
24'b001101010111111000111011, 
24'b111000000110000011011000, 
24'b111111110111111011000111, 
24'b000001100100000110100000, 
24'b000000001101111010011010, 
24'b000001111111001000100001, 
24'b111010100000101110010111, 
24'b000011100111010111100011, 
24'b000001111101101100110000, 
24'b111100001100001100101011, 
24'b000001010001110001010001, 
24'b000000010000010101010100, 
24'b000000100101101100100111, 
24'b111111100100000111100011, 
24'b111111101110000010000110, 
24'b111101110100111101001110, 
24'b000110100000000001110000, 
24'b111001000001111001100111, 
24'b000011011011001100001101, 
24'b111110011001110101010010, 
24'b000011001110000010110110, 
24'b111100010000000010011111, 
24'b000001011010111111001011, 
24'b000000011100111100110000, 
24'b111110011000000010110010, 
24'b000110001101000011111101, 
24'b110011111000110100000011, 
24'b001010010000001101111001, 
24'b000001000111111001000010, 
24'b110101011000111100011111, 
24'b001001011101001000110101, 
24'b111100100000111001011110, 
24'b000010010110000010011111, 
24'b111011100000111101110110, 
24'b0_00011100110000011011010, 
24'b000011011101111011100100, 
24'b111010000000000010001110, 
24'b001000110100000000101011, 
24'b110110010100111100110100, 
24'b000111100000000100110010, 
24'b111101000000111010101101, 
24'b111110100000000100100100, 
24'b000011011110111101100001, 
24'b111110010101111111011010, 
24'b111100111000000011101001, 
24'b001000100110111010101011, 
24'b110100000100000100110011, 
24'b001011010101111101100101, 
24'b111001010011111111110011, 
24'b111111100100000001000101, 
24'b000111100111000000110001, 
24'b110011011011111011001111, 
24'b001101111111001001000100, 
24'b110100001100110100001011, 
24'b000111001001001100001110, 
24'b111110011111110101010110, 
24'b111100010001001000000101, 
24'b001000000010111010110010, 
24'b110100100010000010001101, 
24'b001110001110000000101001, 
24'b110000001000111101100101, 
24'b001111010110000001110000, 
24'b110100100010000001111111, 
24'b000100001011111000100000, 
24'b000100101100001011100010, 
24'b110100011101110101011010, 
24'b001100110011000011010111, 
24'b111001000100000111110001, 
24'b111011111001101110010110, 
24'b001111100000010101010011, 
24'b101010000001101110111110, 
24'b010100111011000111101010, 
24'b110010000111000001011110, 
24'b000101110110111010000110, 
24'b111101111110000100111111, 
24'b000100110000111110010111, 
24'b110100001110111111110100, 
24'b010001111100111110111000, 
24'b101101101010000011101101, 
24'b001011110111111100010001, 
24'b111110011010111110110011, 
24'b111001001010001001111010, 
24'b001001000100101110000011, 
24'b111011011101010100110011, 
24'b111100110011101111001101, 
24'b001001000101001000010101, 
24'b110110010110000000000010, 
24'b000101000100111011011100, 
24'b000001011111000100101110, 
24'b111001111111111101001110, 
24'b000110010101000001100010, 
24'b111101000001111101110110, 
24'b111110011111000011100100, 
24'b000100110001111100001011, 
24'b111010010011000010000010, 
24'b000100110010000000101111, 
24'b111101000000111101010111, 
24'b000001000001000010100011, 
24'b000001000111111110111010, 
24'b111100110110000000000010, 
24'b000100011001111111100001, 
24'b111100010111000001111001, 
24'b000000100011111101100001, 
24'b000011101001000000111111, 
24'b111001110111000001111111, 
24'b000100011011111011110101, 
24'b000001110100000011010101, 
24'b110110001110000000101010, 
24'b001110101100111010101000, 
24'b110011001100000111011000, 
24'b000100001011111011010000, 
24'b000111000000111110100011, 
24'b110001011001000111110011, 
24'b001110011101110101000110, 
24'b111000111011001001100011, 
24'b111101100001111010101101, 
24'b000111111011000001000001, 
24'b111010000001000001010101, 
24'b111110100000111110010101, 
24'b001000101101000001011000, 
24'b110101111010111110011111, 
24'b000100010111000001111000, 
24'b000100100011111110101100, 
24'b110110000000111111000011, 
24'b000111010110000100000111, 
24'b000010101000111001111110, 
24'b110010000011000100111011, 
24'b010011011011111111010001, 
24'b110000101110111011100011, 
24'b000011110111000111111000, 
24'b001000001100111000001101, 
24'b110001110000000100101000, 
24'b001100000110111111110000, 
24'b111010111110111100011101, 
24'b111111001111000110001110, 
24'b000000101101110111100101, 
24'b000101001001001010110110, 
24'b110011100101110010111110, 
24'b001111110101001101100111, 
24'b110011001011110100101001, 
24'b000101010011000110011110, 
24'b000010001110111111010011, 
24'b111010001101111100010100, 
24'b000100101110000101101000, 
24'b111110101000111010000111, 
24'b111111000100000110001000, 
24'b000000100110111000101001, 
24'b000001011111001000111011, 
24'b111100111000110111000010, 
24'b000011000000000110001100, 
24'b111110011011111110101111, 
24'b000000011011111100111010, 
24'b111111101000000011111110, 
24'b000000011010111111110101, 
24'b000001100011111001011011, 
24'b111001100010001100110110, 
24'b001100110011110000011100, 
24'b101111000010001101111101, 
24'b001111101110110110010010, 
24'b110111000010000101100011, 
24'b000000001101111100100011, 
24'b000101101001000011100011, 
24'b111010010101111011011011, 
24'b000001001101000101001100, 
24'b000011001001111011000111, 
24'b111101000100000100001101, 
24'b111101011010111100000011, 
24'b001001110110000100100011, 
24'b110010101101111010001000, 
24'b001001101001000111100100, 
24'b111111101011110110101101, 
24'b110110100111001010111000, 
24'b001110001111110100001001, 
24'b110011011111001011101101, 
24'b000111001101110101111000, 
24'b111100101001000111101100, 
24'b000100010010111010001001, 
24'b110110111111000110001001, 
24'b001101010011110111001000, 
24'b110011000010001100100111, 
24'b000111001110110001001100, 
24'b000000110011001101100100, 
24'b111001100110110110111100, 
24'b000110111011000011101101, 
24'b111100010011111111100001, 
24'b000000111001000000110100, 
24'b111101101100111100100011, 
24'b001000100011000101010011, 
24'b101111100000111100010010, 
24'b010101100110111110100101, 
24'b101011010001000111100001, 
24'b001110001101110101000100, 
24'b111010111011001001100010, 
24'b111101001000111100000100, 
24'b000111000111111100111111, 
24'b111000110010001000010010, 
24'b000100010000110101101111, 
24'b000000000110001001011010, 
24'b111011111011111001000011, 
24'b000101110111000011110100, 
24'b111100000010111111111110, 
24'b111110000101111011100010, 
24'b001001110111001001000011, 
24'b110000001001110011110100, 
24'b001111101010001100011100, 
24'b111000011011110110001101, 
24'b111010010001000101110011, 
24'b010010000011111101000110, 
24'b101001000010000010100110, 
24'b010010000111111011011101, 
24'b111001010101000111000111, 
24'b111011110000110111010100, 
24'b001000011000001001000011, 
24'b111011110011110110111000, 
24'b111011111110001001110010, 
24'b001001011100110101011100, 
24'b111000100111001001110110, 
24'b111110100011111001110001, 
24'b001011101111000000011100, 
24'b101110100111000100101100, 
24'b001111111001111010010000, 
24'b110110010101000001100010, 
24'b000100000100000101110011, 
24'b111100111110110100011010, 
24'b000110011101001100000011, 
24'b110101110010111001001110, 
24'b001001110000111111010001, 
24'b111100100011000101101100, 
24'b111010001110111010100110, 
24'b001100100001000001010010, 
24'b110011100110000010011000, 
24'b000101000010111110011000, 
24'b000110000010111011111011, 
24'b110000100111001011011101, 
24'b010011001111110000000110, 
24'b101111000100001110111001, 
24'b001010110011110110010010, 
24'b111100000001000100011011, 
24'b111110101010111101010000, 
24'b000100101001000101010110, 
24'b111001100001110110011010, 
24'b000111011100001011100100, 
24'b111000011110110110111110, 
24'b000110100001000011000001, 
24'b111011011100000011001110, 
24'b000010001110111001100101, 
24'b111111101001000101011100, 
24'b111111011010111110001111, 
24'b000000101110111110001010, 
24'b111111011001000011000101, 
24'b000000101011111110101110, 
24'b111111000110111101010100, 
24'b000001001000000111001110, 
24'b111110101011110101001111, 
24'b000001110110001100001101, 
24'b111100110101110101000010, 
24'b000101010001000111010111, 
24'b111000101111111101010111, 
24'b000111111100111110111100, 
24'b111001100001000001110001, 
24'b000011001110000001000111, 
24'b000000010111111010000000, 
24'b111101100100001001110111, 
24'b000010000100110110001001, 
24'b000000000101000101011111, 
24'b111101111100000001000001, 
24'b000001110110111010001000, 
24'b000001011001000110010010, 
24'b111001010001111101111110, 
24'b001100000000111011101111, 
24'b110001001000001001010001, 
24'b001110010110110101001100, 
24'b110101000100001001001010, 
24'b000110011001111001111000, 
24'b111101100001000011010111, 
24'b000000001100111110101111, 
24'b000000101100111111000011, 
24'b111111000011000011111010, 
24'b000001010000111000111000, 
24'b111110011001001001010010, 
24'b000001011110110110101100, 
24'b111111101100000111101000, 
24'b111110010011111001111111, 
24'b000011100010000110001111, 
24'b111100000101110111100010, 
24'b000010000100001011000011, 
24'b000001100000110100010110, 
24'b111010110011001001010110, 
24'b000111001011111010011110, 
24'b111001100011000011000100, 
24'b000011101000111011111000, 
24'b111111100000001000011001, 
24'b111111000101110010111100, 
24'b111111100111001110111110, 
24'b000011110101110011000101, 
24'b111000010110001000101100, 
24'b001010001100111010010100, 
24'b110101011011000110011011, 
24'b001001011000110101100110, 
24'b111000001100001110011011, 
24'b000111001000110001010101, 
24'b111000010011001001011111, 
24'b001001001100111111011100, 
24'b110101010001110111111100, 
24'b001011011110001100100001, 
24'b110101001010110100110010, 
24'b001000100100000101100111, 
24'b111011010100000001000001, 
24'b111111111100111010100001, 
24'b000100010100000110000110, 
24'b111001101110111100111101, 
24'b000100100100111110000011, 
24'b000000110110000110110001, 
24'b110111101111110110011100, 
24'b001110101110001001011101, 
24'b101110100011111001000010, 
24'b001111011011000100000110, 
24'b110110011101111100101101, 
24'b000010001111000110010101, 
24'b000100000011110011010010, 
24'b111000001101010011101001, 
24'b001000101011101000110101, 
24'b111001010001010100101110, 
24'b000010001011110011001111, 
24'b000100100111000010111101, 
24'b110011101011000100000110, 
24'b010010010110111010010111, 
24'b101100010011000010011110, 
24'b001110110101000001111010, 
24'b111010101101111100000000, 
24'b111011100111000010110101, 
24'b001001000110111111100011, 
24'b111001110110000000000010, 
24'b111101100000111101000010, 
24'b001011010100000111011110, 
24'b110001010101110110011011, 
24'b001010100110000110010010, 
24'b111101110101000001111110, 
24'b111011011011110100111001, 
24'b000101000100001111111111, 
24'b000000100010110010000101, 
24'b111000110000000110010111, 
24'b001001000001000010001010, 
24'b111100110111111000111111, 
24'b111000100100000110011111, 
24'b001111111001111101101111, 
24'b101111110111111101110100, 
24'b000111001010000100100101, 
24'b000110011010111010111011, 
24'b101110110101000101100010, 
24'b010100000110111000100100, 
24'b110000101111001010000010, 
24'b000111010110110101001110, 
24'b111110001101000111001110, 
24'b000001000001000000110001, 
24'b111101000001110101101011, 
24'b000011100011010001001110, 
24'b000000000111101101100010, 
24'b111001000101001110010000, 
24'b001100110100111000001101, 
24'b110010001111000011001011, 
24'b001000111010111101001011, 
24'b111110101110000110000111, 
24'b111011101110110101111111, 
24'b000100100101001011010010, 
24'b111111110010110111101001, 
24'b111011000110000010010100, 
24'b000110100001000011111110, 
24'b111101000001111000010110, 
24'b111100011100000111101001, 
24'b001000101100111011001001, 
24'b110111011111000001101101, 
24'b000010010011111111101010, 
24'b000111010010000001011101, 
24'b110000010000111100001001, 
24'b010011100001000101010100, 
24'b101110011001111011110110, 
24'b001011110100000000100010, 
24'b111010110011000011100010, 
24'b000000010000111010110110, 
24'b000010010110000010100111, 
24'b111100011101000011010100, 
24'b000100110011110110011110, 
24'b111001010100001100010101, 
24'b001000011011110110011000, 
24'b110111110101000010011110, 
24'b000100011111000101101000, 
24'b000010100010110101001100, 
24'b110101001001001011001011, 
24'b010001010110111000010110, 
24'b101100101001000011000010, 
24'b010000001101000000001111, 
24'b110110011011111110010110, 
24'b000010100100000010101001, 
24'b000010001010111011001100, 
24'b111100011011001000010011, 
24'b000010100101110100101011, 
24'b111111001010001011101011, 
24'b111111011111110111011101, 
24'b000001101101000011100101, 
24'b111100001110000000001010, 
24'b000111010000111111100110, 
24'b110100110100111101100011, 
24'b001101101010000101101001, 
24'b110010111000111001111011, 
24'b001001111010000010101000, 
24'b111001101001000011000101, 
24'b000101011001110111111110, 
24'b110111100111001010001111, 
24'b001101110100110101101110, 
24'b101101110111001010100010, 
24'b010010000010110011001010, 
24'b110011001011010000100110, 
24'b000101000011101101000010, 
24'b000001001011010001001000, 
24'b111101010001110101000010, 
24'b111111101101000011101110, 
24'b000101000010000000001010, 
24'b111000010011000001101101, 
24'b000110010101111000101111, 
24'b111110010010001011010111, 
24'b111100100111110110101110, 
24'b000110011101000000011110, 
24'b111001010100001010100011, 
24'b000101010010101111000100, 
24'b111100000111001110010100, 
24'b000011010000111100000011, 
24'b111101001011111000001100, 
24'b000001011101001101101010, 
24'b000001001001110101111010, 
24'b111100000000111111100101, 
24'b000101011111001011001011, 
24'b111011001101110000011001, 
24'b000010100111001011011101, 
24'b111111010100111110001111, 
24'b000000011001111000100001, 
24'b111110011101001011000110, 
24'b000010100000111000010101, 
24'b111110100101111111111011, 
24'b111110000000000111100100, 
24'b000110000010110101001100, 
24'b111000001000001000011011, 
24'b000101101000111110010111, 
24'b000000010101111001010010, 
24'b111000101110001101101100, 
24'b001011110110101110111101, 
24'b110100000111010000000001, 
24'b000111101010110100100101, 
24'b111110100111000101011001, 
24'b111011110111111111011011, 
24'b000111001000111110111111, 
24'b111000110010111111001001, 
24'b000101010011000100100100, 
24'b111101011001111000100110, 
24'b000000001000000111010011, 
24'b000001100001111011111010, 
24'b111110000111111111100001, 
24'b000000111110000100000110, 
24'b000000111011111010101101, 
24'b111101001011000100011011, 
24'b000011100000111101001101, 
24'b111101101111000001100000, 
24'b111111011111111111100100, 
24'b000011010011111110110010, 
24'b111011110001000011111010, 
24'b000010011101111001010000, 
24'b000001011000000111111101, 
24'b111010110011111001110000, 
24'b000110110100000010001111, 
24'b111010101001000001101101, 
24'b000001110101111100111110, 
24'b000001011011000001001010, 
24'b111101111101000010000001, 
24'b111111000111111100100010, 
24'b000110100000000001101011, 
24'b110011011111000001101111, 
24'b010000011110111101001100, 
24'b101111000110111110011011, 
24'b001101110101001010110001, 
24'b110111011011101100000110, 
24'b000010111101010110101101, 
24'b000001011101110000001110, 
24'b111100000011000001100100, 
24'b000100110111001100110000, 
24'b111010110001101100010011, 
24'b000110001111010000010001, 
24'b110111101001111010000010, 
24'b001010111110111100001110, 
24'b110011100100000110100111, 
24'b001011000000111110100000, 
24'b111010001111111001001000, 
24'b111101110011001011101011, 
24'b001010010101110111001000, 
24'b110000100011000000000000, 
24'b001111101001001001000111, 
24'b110100110000110011011110, 
24'b000100110001001000011001, 
24'b000000100111000000000011, 
24'b111101001001111001010010, 
24'b000010000010000110111011, 
24'b111111111001111111101110, 
24'b111111010001110110100110, 
24'b111111101111010000110010, 
24'b000001111111101101101101, 
24'b111101101111001110000001, 
24'b111111101110111001001000, 
24'b000100111001000000101101, 
24'b110111001011000010000001, 
24'b001000111110111111000001, 
24'b111011111000111101100110, 
24'b111011111011000110000110, 
24'b001011101000110111110000, 
24'b110001100010000111110010, 
24'b001010110011111011011110, 
24'b111101111101111111010111, 
24'b111000000101000101111001, 
24'b001111000110110110111100, 
24'b101110110100001000110001, 
24'b001110011100111010101011, 
24'b110111010100000001000111, 
24'b000001111101000000101011, 
24'b000100100111000010010011, 
24'b110101011011110110001010, 
24'b001111010011010011001110, 
24'b101110101101100101100101, 
24'b001110111000011100010100, 
24'b111000101010100111111000, 
24'b111100010110001111100101, 
24'b001110010011111010001011, 
24'b101011100111111101110100, 
24'b010011101110000110100111, 
24'b110010011011111001000000, 
24'b000110000110000011110111, 
24'b111110011011000001100000, 
24'b000001111111111000111101, 
24'b111010010011001010011011, 
24'b001000110100110110011100, 
24'b111000001111000011111101, 
24'b000001111000000100101110, 
24'b000110010110110011010000, 
24'b110010111111010000011001, 
24'b001111010101110010001001, 
24'b110010110100000110100111, 
24'b001000110101000001001100, 
24'b111011000010111010110001, 
24'b000010111111000011011010, 
24'b111101011011000010110010, 
24'b000010011110110110101000, 
24'b111101111101001100011110, 
24'b000001110001110101011110, 
24'b111101011000000101001100, 
24'b000100101010000000001010, 
24'b111001010110111101011111, 
24'b000110110000000001001111, 
24'b111100000100000010000000, 
24'b111111000011111011100101, 
24'b000101011110000100000100, 
24'b111000101100111111010101, 
24'b000101110001111011101100, 
24'b111101110110001001000111, 
24'b111110100010110011011011, 
24'b000011111011001110100101, 
24'b111010010101110000100001, 
24'b001000000000001111101000, 
24'b110100101011110001010101, 
24'b001110001011001100000100, 
24'b110010001010111000011100, 
24'b001000101000000001110001, 
24'b000000100011000011111001, 
24'b110110001101111000001101, 
24'b001110101110001000111101, 
24'b110010110110111000011011, 
24'b000110110111000101000010, 
24'b111111100110111100110010, 
24'b111110001001000011100101, 
24'b111110101000111001110001, 
24'b000111100101001001111110, 
24'b110011110101110011001100, 
24'b001011101010001101010000, 
24'b111010001011110100111101, 
24'b111101011101000111010100, 
24'b001001110000111100010011, 
24'b110010100111000001000011, 
24'b001101100001000001001010, 
24'b110100011111111011100111, 
24'b001000110111001001101001, 
24'b111001111111101111111101, 
24'b000010111100010100110100, 
24'b111111111101101011011010, 
24'b111110101100001101110101, 
24'b111111101011111101101110, 
24'b000101001010110110100100, 
24'b110100101111010000001110, 
24'b001111100101110000011101, 
24'b110000100001001000110111, 
24'b001010110101111111010000, 
24'b111100000000111011111110, 
24'b111110010110000011011101, 
24'b000011111010000000110011, 
24'b111101000111111011001010, 
24'b000000100110000101011110, 
24'b000000110010111101101100, 
24'b111111100011111101101001, 
24'b111111000110000101100011, 
24'b000010000101111010001000, 
24'b111101011111000100010111, 
24'b000010011110111100110010, 
24'b111101101001000011101001, 
24'b000001110111111011011011, 
24'b000000000000000011100011, 
24'b111100001001000001001101, 
24'b001000110000110111010000, 
24'b110011101111001111011101, 
24'b001100000001101110101110, 
24'b111000001110001100101010, 
24'b000010001011111100001011, 
24'b000000101101111011110110, 
24'b000001101100000110100101, 
24'b110111110111111101111110, 
24'b001110000101111001010100, 
24'b110001101000001110011010, 
24'b000111001001101111010101, 
24'b000100100001001100010110, 
24'b110001110000111100000100, 
24'b010000100101111011110001, 
24'b110101011110001000110011, 
24'b000000011010110110111110, 
24'b000111001110000110111010, 
24'b111000010011111010101000, 
24'b000001010101000110100001, 
24'b000111011001110101101101, 
24'b110011001001001110110100, 
24'b001100001001101110100101, 
24'b111001101011010000000110, 
24'b111111001111110101100101, 
24'b000101100010000001101011, 
24'b111001010111000111101101, 
24'b000101000111110000111011, 
24'b111101011011010010110001, 
24'b111111111000101101011111, 
24'b000011001100001111100110, 
24'b111001010001110100000101, 
24'b001001101010001001000001, 
24'b110110000111111000110010, 
24'b000101111110000101100111, 
24'b000001001101111100111100, 
24'b110111101001111111001000, 
24'b001011101010000101010011, 
24'b110110100111110111101000, 
24'b000011011100001000100011, 
24'b000001110100111010011100, 
24'b111101100011000000101010, 
24'b111101101011000100001010, 
24'b001001101001111000100101, 
24'b110001000100001000110100, 
24'b001111010101110111000000, 
24'b110100101101001000101100, 
24'b000110001010111000001001, 
24'b111100101110000101111001, 
24'b000011101111111101100101, 
24'b111010001111111110010001, 
24'b000110101011000100100111, 
24'b111010110000111011111000, 
24'b000010110111111111101010, 
24'b111101101101000111001010, 
24'b000101001111110010111111, 
24'b110101101000001110101101, 
24'b001110000101110101000000, 
24'b110010111111000011100010, 
24'b000110110111000100000110, 
24'b000001000000110111101010, 
24'b111010011100000111101110, 
24'b000011101001111100100111, 
24'b000011110111111110010111, 
24'b110011101101000100010011, 
24'b010000100100111100110011, 
24'b110001100000111111001011, 
24'b001000011100000101011001, 
24'b111100100000111000000111, 
24'b000100000010000111001010, 
24'b110101011011111100001100, 
24'b010011011100111111111111, 
24'b100110111011000010000110, 
24'b010111110101111110100101, 
24'b101111110111111110110010, 
24'b000110001111000011101000, 
24'b000000101010111100010110, 
24'b111110100001000000100000, 
24'b111100111110000100110011, 
24'b001001010111110110001011, 
24'b110010100010001100011110, 
24'b001101010100110011110010, 
24'b110110011000001010010010, 
24'b000100110000110111010111, 
24'b111111001000001000011001, 
24'b111110101000110111001000, 
24'b000010110111001000010010, 
24'b111011001110111010110100, 
24'b000111010110000000000111, 
24'b110110100111000100100001, 
24'b001001010100111001111111, 
24'b111001100110000011100100, 
24'b000001101100000000110011, 
24'b000010010101111100100111, 
24'b111100110101000001011010, 
24'b000000010000000100110000, 
24'b000100100100110100100000, 
24'b111000010110001110011010, 
24'b000101111101110100110100, 
24'b000001001011000011100001, 
24'b110100111101000100000110, 
24'b010010111110111000100100, 
24'b101011001101000101100011, 
24'b001111010110111110101011, 
24'b111010111100111111010000, 
24'b111010100111111101111101, 
24'b001011110001001000101011, 
24'b110011100000110001001010, 
24'b001001001001010000010000, 
24'b111011010000110100100110, 
24'b000001100101000010101100, 
24'b000000011001000101010110, 
24'b111101001101110111001101, 
24'b000111000000000110100100, 
24'b110011100111111111011101, 
24'b010000001110111001110000, 
24'b110000100001001011011010, 
24'b001001011101110001111110, 
24'b111111011001001110000111, 
24'b111001011011110100001100, 
24'b001000110011000111001011, 
24'b111001110101111111001100, 
24'b000010011010111010100101, 
24'b111110000100001000111000, 
24'b000110011111111000100001, 
24'b110010110000000001011001, 
24'b010000101110000110101100, 
24'b110011100010110011010010, 
24'b000000110011001101101100, 
24'b001100111111110110101101, 
24'b101010010101000001101110, 
24'b010100110001000101111111, 
24'b110100100010110100010001, 
24'b111111100000001111001010, 
24'b001000111010101111001110, 
24'b110100110000010000101101, 
24'b001001110101110001101110, 
24'b110110101111001000111101, 
24'b001100011100111110010100, 
24'b101110000100111011001111, 
24'b010101000011000111000101, 
24'b101110010000111100010000, 
24'b001000000101111100100011, 
24'b000011010010001010010010, 
24'b110101101101110011010111, 
24'b001001110010001001010110, 
24'b111100011101111101000101, 
24'b111100111001111101110110, 
24'b000101100011000010101000, 
24'b111100111110000001010100, 
24'b111110111011111001100010, 
24'b000010100011001000111100, 
24'b000000000011111001000010, 
24'b111011111010000001101101, 
24'b000101001010000011111110, 
24'b111110111100111000010010, 
24'b111010000001001001010010, 
24'b001010101011110110001101, 
24'b110111010100001010010011, 
24'b000000011001110101100100, 
24'b001001000101001000111001, 
24'b110010100111111011000000, 
24'b001001101111111111111011, 
24'b111111000000000011100011, 
24'b111001101100111100111000, 
24'b000110111001111110111101, 
24'b111111100010000110000110, 
24'b110111101101110111101010, 
24'b001101100000000101111110, 
24'b110011100001111111011011, 
24'b000111101010111100000100, 
24'b111100001000000100001111, 
24'b000100010101111111110111, 
24'b111000010110111010110011, 
24'b001001000111000111100011, 
24'b111011001110111011010011, 
24'b111011010001111110001011, 
24'b001110000111001000000111, 
24'b101111000100110101011100, 
24'b001010101011001000100110, 
24'b000001001001111011001010, 
24'b110100110011000011000000, 
24'b001101100010111011000101, 
24'b111000010111001001001011, 
24'b111110101011110100000000, 
24'b000110100010001001111001, 
24'b111011100011111110000010, 
24'b111101001011110110101001, 
24'b001001100101010011111001, 
24'b110101001011100110001110, 
24'b000101111001011001011000, 
24'b000001011111101100011111, 
24'b111001101000001010110101, 
24'b000110011011111101100010, 
24'b111100111001111101000100, 
24'b000000001101000011111010, 
24'b111111110000111111001101, 
24'b000010110101111011101100, 
24'b111010110110001000010010, 
24'b000100110000110111110110, 
24'b111110011001000010111111, 
24'b111110001011000101011000, 
24'b000010110010110010111000, 
24'b111111011010010000100001, 
24'b111101010000110001101010, 
24'b000100001000001000101011, 
24'b111110001010111100100000, 
24'b111100110110000010000001, 
24'b001000001000111011101000, 
24'b110101010011000111100101, 
24'b001010100011111000010011, 
24'b110110110110000010111011, 
24'b001000001101000101001000, 
24'b111000001100110011110100, 
24'b000110100000001110011001, 
24'b111101010111110101011001, 
24'b111100001011000011001000, 
24'b001010110110000100010000, 
24'b110000011101110111001010, 
24'b010000010001001010100101, 
24'b110010010001110100110001, 
24'b001010010011001100100001, 
24'b110111111011110001111101, 
24'b000111011101001101101001, 
24'b111001000101110110111010, 
24'b000100110100000000011101, 
24'b111111010010001001010100, 
24'b111100000110110000010010, 
24'b000110111110001111100000, 
24'b111000100000110111001100, 
24'b000110011010111111001010, 
24'b111010000110001000100101, 
24'b000111110011110101000101, 
24'b110011111111000111100100, 
24'b010000100101111110111111, 
24'b101101000010111010110110, 
24'b010001100100001000011001, 
24'b110011011000110111110111, 
24'b000101111010000101011111, 
24'b000000010011111101111000, 
24'b111011111010111111010001, 
24'b000100011110000010100011, 
24'b111110100110111100111101, 
24'b111011111000000010001010, 
24'b001010001101000000001011, 
24'b110001100111111100100010, 
24'b001110101111000110100100, 
24'b110100111100111000000111, 
24'b000101000110000110010100, 
24'b000000001101111110001100, 
24'b111101011001111011110110, 
24'b000010000110001001100000, 
24'b111111010011110011101000, 
24'b000000110101001100010011, 
24'b111101000100110101110101, 
24'b000100111001000111110110, 
24'b111100011111111001010000, 
24'b111101011010000111001101, 
24'b001011001110110111110011, 
24'b101110100010001000010010, 
24'b010001000011111001100110, 
24'b110110010000000010101101, 
24'b000000010101000001101010, 
24'b000100100000111010110101, 
24'b111111010110000111000000, 
24'b110110000110111000101000, 
24'b010100010111000111001011, 
24'b101000110111111000111011, 
24'b001111010110000110111100, 
24'b111111100111111010010000, 
24'b110001111000000010100101, 
24'b010101101000000010011110, 
24'b101011100010111000001100, 
24'b001110010100001011000000, 
24'b110111001110110101111111, 
24'b000111001010000100101100, 
24'b110111011100000011000011, 
24'b001001011100110110000000, 
24'b111001000011001101001011, 
24'b000001011111110100101111, 
24'b000011110101000101000010, 
24'b111010011000000011010111, 
24'b000010111100110100110000, 
24'b000010011011010000100011, 
24'b111000100010101101111011, 
24'b001010010110001111100111, 
24'b110100111001110110010000, 
24'b001010100110000001110100, 
24'b110111001100000110001110, 
24'b000100101010110011100111, 
24'b000010100111001111100101, 
24'b110100100011110000000110, 
24'b010001111011001110111010, 
24'b101110001011110001101000, 
24'b001010001001001111001101, 
24'b000001010011101111010010, 
24'b110110011100010001000000, 
24'b001001000111110001101100, 
24'b000000010010001000100010, 
24'b110011000001111110101000, 
24'b010101010100111011100001, 
24'b101011011001000111000111, 
24'b001100011011111001100001, 
24'b111101000101000100011001, 
24'b111110000011111100110011, 
24'b000000110110000100001011, 
24'b000010010101111001001000, 
24'b111110000000001001100010, 
24'b111011110111110101101011, 
24'b001100101111001000011111, 
24'b101110111100111011100010, 
24'b001100001100111111100101, 
24'b000000110110000100110011, 
24'b110000111010111000011001, 
24'b010110001110001000000010, 
24'b101110000010111010010100, 
24'b000101000000000000110001, 
24'b001001001101000101100001, 
24'b101110100111110100111110, 
24'b010000111100001101011001, 
24'b110101011011110100110000, 
24'b000011100011000101010011, 
24'b000000101000000001110111, 
24'b111101111101111000111110, 
24'b000011010001000111111100, 
24'b111001110001111011100000, 
24'b001010001010111110011001, 
24'b110100000000000111111101, 
24'b001001001000110011010001, 
24'b111110001010001111010000, 
24'b111001110000110000011000, 
24'b001010101001001110011010, 
24'b110111000110110011110000, 
24'b000010011001001010001010, 
24'b000100110111110110100001, 
24'b110111010000001011001111, 
24'b000111101001110000110110, 
24'b111100111010010011001110, 
24'b111110011011101011101001, 
24'b000011011100010000011111, 
24'b111110011011110111101001, 
24'b111101000100111111110010, 
24'b000111110101000100011000, 
24'b110101000101111110100110, 
24'b001010110101111000110001, 
24'b111000100001010000011011, 
24'b000010000100101011010110, 
24'b000011000010010001100011, 
24'b111010110001110110101001, 
24'b000010111000000001001111, 
24'b000011011011000010100100, 
24'b110101011111111110100010, 
24'b001110001110111110101100, 
24'b110100011011000001101011, 
24'b000011001001000001111001, 
24'b000111000010111000110101, 
24'b110010011011001010000001, 
24'b001101001000111000000001, 
24'b111001100101000010100000, 
24'b111101110110000010001001, 
24'b000111100100111101101110, 
24'b111000101110111110000000, 
24'b000010111100000110100001, 
24'b000001010100111001110011, 
24'b111110000110111111010000, 
24'b111110011110001010110000, 
24'b000110000100101111001010, 
24'b111000010100001101100101, 
24'b000100011010111110111000, 
24'b000010011010110001100100, 
24'b110111000101011000101110, 
24'b001011011001100111011101, 
24'b110111100100001111001000, 
24'b000001100010111101001001, 
24'b000110010101111010111110, 
24'b110011100001000101000110, 
24'b001111111101000000101010, 
24'b101110111011111001000000, 
24'b010000100111001001011110, 
24'b110000111011111000110011, 
24'b001100110010000010111001, 
24'b110101110000111111110100, 
24'b001000010110000000110000, 
24'b111000011010111100100010, 
24'b000111100001000101100110, 
24'b111001100001111010110011, 
24'b000010110111000010100000, 
24'b000011101001000000101000, 
24'b110100111011111101110010, 
24'b010000001001000001110000, 
24'b101111110001111111110110, 
24'b001011010000111110110111, 
24'b111100000101000001011110, 
24'b111110000100111110111100, 
24'b000011111100000000011101, 
24'b111101011100000000010000, 
24'b000000100110111110100010, 
24'b111111001000000011010111, 
24'b000100000001111010110100, 
24'b111000001000000101010111, 
24'b001001010110111101001101, 
24'b111001011101111110000001, 
24'b000000100001000110011101, 
24'b000101100110111000100000, 
24'b110111011001000011101001, 
24'b000111011000000011101000, 
24'b111100101011110101101100, 
24'b111111000000001100011101, 
24'b000011111011110111010100, 
24'b111010011110000001010110, 
24'b000111001000000100110001, 
24'b110110101001111010100010, 
24'b001011001110111111111100, 
24'b110101010011001000101101, 
24'b000110100100110000110010, 
24'b111111111011001111100010, 
24'b111010110110110110111000, 
24'b000101010010111111011100, 
24'b000000111110001000011010, 
24'b110101000010110101011101, 
24'b010011010100000110100101, 
24'b101010111111000000011110, 
24'b001110101100111001110110, 
24'b111100101000000111010100, 
24'b111000111001111100010100, 
24'b001011101110111101110000, 
24'b110110111111000111000100, 
24'b000001100010110111100101, 
24'b000110001100000110010010, 
24'b110101100001111101011110, 
24'b001010011101111111100000, 
24'b111000000110000001100001, 
24'b000101011011111111001100, 
24'b111011011000111111100101, 
24'b000101001110000001001000, 
24'b111010001100111110101100, 
24'b000101010011000001101110, 
24'b111100011101111101000001, 
24'b000001011111000100110011, 
24'b000000000101111010001110, 
24'b111110111001000100100010, 
24'b000010010100111111010110, 
24'b111011101101111011011111, 
24'b000110111001001000101010, 
24'b110111000110110110010010, 
24'b001001001011000111001101, 
24'b111000100110111101100010, 
24'b000100101101111101110111, 
24'b1_11101000100000100101010, 
24'b111100000111111010100011, 
24'b000111001000000111110010, 
24'b110101100111110111010111, 
24'b001101001100000111111010, 
24'b110000111110111010010001, 
24'b001111100101000010011100, 
24'b110001011011000001011101, 
24'b001100000011111010100101, 
24'b110111101111001000111010, 
24'b000011101011110100100100, 
24'b000001001000001100101110, 
24'b111010100011110011010011, 
24'b001000110001001011011101, 
24'b110101011011110110110010, 
24'b001010101010000110010110, 
24'b110110111110111100101111, 
24'b000101111100000000010100, 
24'b111110001010000010001100, 
24'b111101010110111011111100, 
24'b000110111101000101010000, 
24'b110101100010111010010001, 
24'b001100101110000101101011, 
24'b110010100100111010110100, 
24'b001100100010000100011011, 
24'b110101111000111100011101, 
24'b000110100011000010101110, 
24'b111101110001111110000010, 
24'b111101110001000001011010, 
24'b000110011000111110111010, 
24'b110110011001000001000001, 
24'b001011100100111110101101, 
24'b110100000011000001111000, 
24'b001010101101111101001011, 
24'b111000000100000100000100, 
24'b000011111100111010011010, 
24'b000000101111000111010010, 
24'b111010011111110111000001, 
24'b001001110000001010100001, 
24'b110011001101110100010000, 
24'b001110001100001100011111, 
24'b110010011010110011011001, 
24'b001011000000001100000100, 
24'b111001011000110101001011, 
24'b000000111101001000111111, 
24'b000101010011111001010111, 
24'b110100101110000011111111, 
24'b010000010000111110110100, 
24'b101100011111111110011110, 
24'b010100101010000100000100, 
24'b101100011011111001110100, 
24'b010000100011000111110010, 
24'b110011111010110111001110, 
24'b000111000000001001000110, 
24'b111101111001110111010001, 
24'b111110010000000111101010, 
24'b000100000100111010000011, 
24'b111011100011000011110001, 
24'b000011000111111110101100, 
24'b111111100110111110110100, 
24'b111101000100000011011100, 
24'b000110000101111010110111, 
24'b110111110011000110000010, 
24'b001000110001111010000011, 
24'b111000100111000100111011, 
24'b000100001111111101000000, 
24'b000000010001000000011111, 
24'b111010101001000010001111, 
24'b001010000101111011010101, 
24'b110010011110000110011000, 
24'b001111000001111001000100, 
24'b110001110111000110001010, 
24'b001010110110111011111111, 
24'b111010011000000000110101, 
24'b111111001000000011000000, 
24'b000111101010111001001100, 
24'b110010001010001010000000, 
24'b010010100110110100000101, 
24'b101010100110001100001100, 
24'b010110001100110101010110, 
24'b101010110111000111011011, 
24'b010010110111111101000010, 
24'b101111111110111101111100, 
24'b001101011101000110111101, 
24'b110100010101110101000110, 
24'b001011000110001101010100, 
24'b110100010011110010001000, 
24'b001101001010001100100010, 
24'b110001000101110110011111, 
24'b010000010010000101011010, 
24'b101111011010111111001101, 
24'b001111011011111100011000, 
24'b110011011001000111010101, 
24'b001000010011110110000101, 
24'b111100111100001011011001, 
24'b111101100111110100001000, 
24'b000111001101001011110010, 
24'b110101010110110100011111, 
24'b001100001100001011100001, 
24'b110100011011110011111100, 
24'b001001000000001101010010, 
24'b111011000010110001000100, 
24'b000000001100010000101001, 
24'b000100100000101110000100, 
24'b110111101111010010010011, 
24'b001010100101101110101110, 
24'b110100110111001110110011, 
24'b001010000101110101000110, 
24'b111000010010000110000010, 
24'b000100101101111111001011, 
24'b111110010000111100000010, 
24'b111111011110000111101001, 
24'b000001101010110110011001, 
24'b111110100100001001100101, 
24'b111111111110111000010111, 
24'b000010010100000100001001, 
24'b111011000111000000010001, 
24'b000111001010111011001010, 
24'b110111011100001000110010, 
24'b001000101111110100011110, 
24'b111000011010001100101011, 
24'b000101010000110011101111, 
24'b111101111001001010100100, 
24'b111110101101110111111001, 
24'b000100011111000101100000, 
24'b111001000100111100101000, 
24'b001000011001000010001100, 
24'b110111001110111101110111, 
24'b001000001110000011001100, 
24'b111000111100111011000100, 
24'b000101101100000110111101, 
24'b111011100000110111010111, 
24'b000011110100001001100010, 
24'b111100001111110110101101, 
24'b000100010101000111111001, 
24'b111010101110111010011111, 
24'b000110010010000010100101, 
24'b111001000001000000010111, 
24'b000111000101111101001011, 
24'b111001100110000100010101, 
24'b000100111011111011010010, 
24'b111101001101000011111111, 
24'b000000010111111101100100, 
24'b000010000000000000011111, 
24'b111100000101000001011001, 
24'b000101000100111101010011, 
24'b111010101101000011001010, 
24'b000100101011111101010010, 
24'b111100101001000001100001, 
24'b000001110000000000001001, 
24'b111111110100111110010000, 
24'b111111000110000010111001, 
24'b000001001110111100110001, 
24'b111111011011000010101010, 
24'b111111000000111110110001, 
24'b000011010101111111011000, 
24'b111001110110000010100011, 
24'b001001000110111100000010, 
24'b110100001011000100011101, 
24'b001110000010111100010010, 
24'b110000011011000001110101, 
24'b010000010110000000111110, 
24'b101111101010111011110000, 
24'b001111101110000111011001, 
24'b110001011110110110001100, 
24'b001100111000001011000001, 
24'b110101001011110101001000, 
24'b001000010110001001011001, 
24'b111010100011111001000100, 
24'b000010000011000100000100, 
24'b000001110011111110100001, 
24'b111001111111111111110000, 
24'b001010010100000000101100, 
24'b110001100011000000010111, 
24'b010001111111111101001110, 
24'b101011100010000110000111, 
24'b010101011111110110001110, 
24'b101011001000001101000111, 
24'b010010100011110000100010, 
24'b110001010111010000100000, 
24'b001001101001101111111100, 
24'b111011111010001110010100, 
24'b111110101101110100010011, 
24'b000101110110001000110010, 
24'b110111000101111001110011, 
24'b001010010000000100011111, 
24'b110110010100111100001000, 
24'b000111011100000100011011, 
24'b111011111110111010000111, 
24'b000000000110000111110010, 
24'b000011101000110110011100, 
24'b111001100011001010101000, 
24'b000111111001110101011000, 
24'b111000010110001001010111, 
24'b000101111001111001000001, 
24'b111101000101000011110011, 
24'b111111010110111111101001, 
24'b000100000110111101001110, 
24'b111001010100000101000101, 
24'b000111110101111001101110, 
24'b111000110110000110010010, 
24'b000100100110111010101001, 
24'b111111100010000011111011, 
24'b111011010000111101011101, 
24'b001010010011000001110000, 
24'b110000101000111110000010, 
24'b010011001110000011011000, 
24'b101010101110111010001001, 
24'b010101010001001001000011, 
24'b101100110101110011100111, 
24'b001111010010001111001101, 
24'b110101110010101111000011, 
24'b000100100110010001001011, 
24'b000000110110110000001111, 
24'b111010100010001100111000, 
24'b001000110111110111000110, 
24'b110101001110000100100000, 
24'b001011010111111111101101, 
24'b110101001010111100111001, 
24'b001001101111000101010011, 
24'b110111100001111001110011, 
24'b000111101001000101111001, 
24'b111000100000111011001100, 
24'b001000001011000011011111, 
24'b110110011001111101100110, 
24'b001011100100000010000011, 
24'b110010011110111101011001, 
24'b001111000101000100000110, 
24'b110000010001111001110100, 
24'b001111001010001000011011, 
24'b110010110010110101101101, 
24'b001010000000001011010010, 
24'b111010001101110100111101, 
24'b000001001000001001100010, 
24'b000011011101111001001001, 
24'b111000101010000011011101, 
24'b001010000101000000000101, 
24'b110100101110111100110111, 
24'b001010111010000101001111, 
24'b110110111011111010000001, 
24'b000110001010000101010101, 
24'b111101010110111100100000, 
24'b111111001000000000111010, 
24'b000011111000000001111001, 
24'b111010000110111011101110, 
24'b000110110001000101110001, 
24'b111001100110111001111111, 
24'b000100111110000100111111, 
24'b111101001101111101000101, 
24'b000000011001000000001100, 
24'b000001111000000010101011, 
24'b111100011101111010111001, 
24'b000100011101000110101100, 
24'b111011100000111000110011, 
24'b000011110100000110100100, 
24'b111101010010111010111110, 
24'b000001100100000010111110, 
24'b111111001110111111001110, 
24'b000000101101111110111011, 
24'b111110011001000010001111, 
24'b000011011101111101011110, 
24'b111001110110000010000011, 
24'b001001010110111111000110, 
24'b110011011001111111011110, 
24'b001111011010000001111110, 
24'b101110101110111100111100, 
24'b010001111000000011101000, 
24'b101110111011111100011011, 
24'b001110110111000011000001, 
24'b110100011100111101111010, 
24'b000111100011000001000110, 
24'b111100101001111111101111, 
24'b111111100110111111101101, 
24'b000011010010000000011111, 
24'b111011000010111111100111, 
24'b000101010000000000001000, 
24'b111011110001000000000011, 
24'b000010001111000000000000, 
24'b000000010100111111100100, 
24'b111101000100000001001111, 
24'b000101000101111101110001, 
24'b111001101010000011001111, 
24'b000110011110111100000100, 
24'b111010100110000100000010, 
24'b000011010101111100101110, 
24'b111111011100000001100111, 
24'b111101100100000000111101, 
24'b000101001001111011110111, 
24'b111000111001000111100100, 
24'b000111111101110101001010, 
24'b111000011001001101100110, 
24'b000110000100110000100010, 
24'b111100011101010000010101, 
24'b000000011111101111110101, 
24'b000010101011001111001111, 
24'b111010100000110010001111, 
24'b000111100111001100001011, 
24'b110111001110110101010000, 
24'b001000111101001001101111, 
24'b110111101010110110110010, 
24'b000111001110001001000011, 
24'b111001111111110110111101, 
24'b000101000111001000111000, 
24'b111011001001110111110101, 
24'b000101011110000110101011, 
24'b111001000011111011110011, 
24'b001001001000000000111000, 
24'b110100011000000011000111, 
24'b001110000100111000101010, 
24'b110000000100001011011001, 
24'b010000111001110001010101, 
24'b101111010100010000110110, 
24'b001111011000101110011101, 
24'b110010111010010000110001, 
24'b001010010000110001011010, 
24'b111000101101001011010110, 
24'b000100110100111000100100, 
24'b111100110100000011011000, 
24'b000010101101000000011001, 
24'b111100101011111100100100, 
24'b000100110111000101100000, 
24'b111001001001111001100010, 
24'b001000101100000110010110, 
24'b110110010001111010110000, 
24'b001001011110000011011010, 
24'b111000011111111111000000, 
24'b000011110110111110010000, 
24'b000001010011000100101011, 
24'b111000101101111000011010, 
24'b001101011111001010010111, 
24'b101101000101110011001010, 
24'b010110111001001110111011, 
24'b100111001101101111100011, 
24'b011000010100010001010010, 
24'b101010011011101110101101, 
24'b010001000010010000011011, 
24'b110100100111110001010111, 
24'b000101100101001100000100, 
24'b111111011111110111001000, 
24'b111101000000000101010101, 
24'b000100011101111110001101, 
24'b111100010011111110100111, 
24'b000000111110000011111100, 
24'b000011001010111010011000, 
24'b111000000011000110010110, 
24'b001100011101111001110011, 
24'b110000001001000101010111, 
24'b010001100011111011111010, 
24'b101110110010000010101110, 
24'b001110111001111110100001, 
24'b110101000101000000101010, 
24'b000101111100111111101111, 
24'b111111010100000000010001, 
24'b111011111001111111100010, 
24'b000111110010000000101010, 
24'b110110000011111111011011, 
24'b001010011111000000000010, 
24'b110110011011000001000110, 
24'b000111100111111101010011, 
24'b111010111001000100101000, 
24'b000010101010111001011100, 
24'b111111010011001000001010, 
24'b111111101010110110111011, 
24'b000000010111001001000101, 
24'b000000100101110111111011, 
24'b111101101100000110001010, 
24'b000100100000111100011101, 
24'b111001001110000000101101, 
24'b001000111000000001111101, 
24'b110101011100111100000100, 
24'b001011101111000100111100, 
24'b110011101001111011010000, 
24'b001100100101000011011000, 
24'b110011100001111110111010, 
24'b001100001100111110010001, 
24'b110100001101000100101001, 
24'b001011010100111000111000, 
24'b110101010001001000110010, 
24'b001010000010110110101010, 
24'b110110110101001000110001, 
24'b001000001011111000110110, 
24'b111000111000000100110011, 
24'b000110001111111101111001, 
24'b111010010111111111011111, 
24'b000101101001000010101101, 
24'b111001101011111011110011, 
24'b000111110111000100111111, 
24'b110101111010111010111001, 
24'b001100111011000100110011, 
24'b110000000110111011101110, 
24'b010010101100000011111000, 
24'b101011001110111100010000, 
24'b010101110110000011111110, 
24'b101010011000111011100110, 
24'b010100000001000100111001, 
24'b101110110101111010111110, 
24'b001101011100000100100010, 
24'b110110110010111100111100, 
24'b000101000010000000011110, 
24'b111110101001000011001110, 
24'b111110100110111000010010, 
24'b000011001001001100101000, 
24'b111100001111101110101010, 
24'b000011011111010101010001, 
24'b111101011110101000001100, 
24'b000001010001011000100010, 
24'b111111111101101000110011, 
24'b111111000101010011111000, 
24'b000001100001110001001001, 
24'b111110001110001000101010, 
24'b000001110110111110000010, 
24'b111110000101111011011110, 
24'b000010001111001010001000, 
24'b111101000000110001101000, 
24'b000100001100010000111111, 
24'b111010001100101110001001, 
24'b000111101001010001001110, 
24'b110110100101110000100101, 
24'b001010110101001100111110, 
24'b110100011000110101101100, 
24'b001011100111000111111101, 
24'b110101010000111001110110, 
24'b001001001001000101001001, 
24'b111001000001111011001100, 
24'b000100100011000101000101, 
24'b111101110111111010010101, 
24'b000000000000000110010011, 
24'b000001110000111001010111, 
24'b111100111100000110100000, 
24'b000100000100111010001100, 
24'b111011000111000100100110, 
24'b000101101100111101000100, 
24'b111001011010000001000110, 
24'b000111101010000000101101, 
24'b110111001100111101110001, 
24'b001001110100000011010100, 
24'b110101100111111100001101, 
24'b001010001110000011101011, 
24'b110110111101111101000000, 
24'b000110110010000001111000, 
24'b111100100110111111100001, 
24'b111111001000111111000011, 
24'b000101101001000010010100, 
24'b110101100100111100100100, 
24'b001110101110000100000111, 
24'b101110000000111011110000, 
24'b010100000001000011110100, 
24'b101011011000111101010000, 
24'b010011111101000001000000, 
24'b101101101101000001010111, 
24'b010000001000111011110000, 
24'b110010000100000111100011, 
24'b001100001011110101000000, 
24'b110100110101001110010111, 
24'b001011000011101110101101, 
24'b110100010001010011011111, 
24'b001100111100101011011000, 
24'b110001110000010100100001, 
24'b001111001111101100111110, 
24'b110000100010010000001111, 
24'b001110101000110011100111, 
24'b110011011000000111110101, 
24'b001001100100111100111010, 
24'b111010010010111110101100, 
24'b000001011101000100111011, 
24'b000010101110111000101101, 
24'b111001100011001000010011, 
24'b001001010110111000000001, 
24'b110100110001000110101000, 
24'b001100000111111011010010, 
24'b110011111001000010110110, 
24'b001011011100111110010101, 
24'b110101101001000001101101, 
24'b001001000110111100110001, 
24'b111000000111000110010011, 
24'b000110110001110101011011, 
24'b111010001111001111100001, 
24'b000100110110101011101101, 
24'b111100000111010111111111, 
24'b000010111001100110001010, 
24'b111110010001011001001100, 
24'b000000100100101010010000, 
24'b000000100100001111101100, 
24'b111110100100111000011100, 
24'b000001111001111110010011, 
24'b111110001101001010111011, 
24'b000001000101101101000110, 
24'b000000010000011000011110, 
24'b111110000000100101001001, 
24'b000011111110011001101001, 
24'b111010001010101011000010, 
24'b000111010011001101011100, 
24'b110111111000111011111010, 
24'b001000000111111010001111, 
24'b111000110110001110110011, 
24'b000101010101101010001110, 
24'b111101010000011001110011, 
24'b111111101001100101100111, 
24'b000011110001010111101010, 
24'b111000101110101101111110, 
24'b001010100101001010011110, 
24'b110010011011111101111001, 
24'b010000001000111010001010, 
24'b101101111000001100010111, 
24'b010011011111101111011000, 
24'b101011110101010010010001, 
24'b010100000110101110101101, 
24'b101100110011001110000100, 
24'b010001011100110110110000, 
24'b110001001100000011101010, 
24'b001011011111000001111110, 
24'b111000011100111001000110, 
24'b000011010111001010101111, 
24'b000000110010110010110001, 
24'b111011011110001110100000, 
24'b000111100000110001010010, 
24'b110110100100001110010101, 
24'b001010010000110010010110, 
24'b110110000101001101000011, 
24'b001000101101110011011011, 
24'b111001000011001100010111, 
24'b000101000101110011110001, 
24'b111100011011001011111110, 
24'b000010110011110100100111, 
24'b111101000000001010010000, 
24'b000100001010110111100010, 
24'b111001111000000110001100, 
24'b001000100011111100011101, 
24'b110101000101000000111010, 
24'b001100101010000001011101, 
24'b110010101100111100110100, 
24'b001100100010000100000110, 
24'b110101110000111011111001, 
24'b000110100011000011010111, 
24'b111110001101111101111100, 
24'b111100100100000000101000, 
24'b001000011110000000100101, 
24'b110011010011111110101111, 
24'b001111100011000001001111, 
24'b101111010100111111100010, 
24'b001111111101111111000110, 
24'b110010100000000010100010, 
24'b001001101101111011111110, 
24'b111010111011000101000001, 
24'b000000001110111010111100, 
24'b000100010000000100000110, 
24'b111000001001111101111100, 
24'b001010001011111111010001, 
24'b110100111111000011111001, 
24'b001010011100111001001001, 
24'b110111011100001001000110, 
24'b000101110001110101111011, 
24'b111101100111001001011111, 
24'b111110111011111000110000, 
24'b000100001111000011100010, 
24'b111001010100000001010100, 
24'b001000010000111001010100, 
24'b110111010001001011111110, 
24'b001000001000101111100000, 
24'b111001011111010011110011, 
24'b000100001001101010011110, 
24'b111110101111010101100100, 
24'b111110010001101011111101, 
24'b000100011111010001010011, 
24'b111001010101110010010000, 
24'b000111111101001001110111, 
24'b110111110000111001111001, 
24'b000111100001000010110110, 
24'b111010000111111111101100, 
24'b000011101000111110100100, 
24'b111110110101000010011001, 
24'b111110111010111101011000, 
24'b000010101101000010010111, 
24'b111100101100111110010110, 
24'b000010110011000000100111, 
24'b111110111000000000101111, 
24'b111110100011111101101011, 
24'b000100100101000100010010, 
24'b111000010010111001011101, 
24'b001010010100001001000011, 
24'b110100000010110100010101, 
24'b001100010100001110001111, 
24'b110100101100101111100011, 
24'b001001000110010010000110, 
24'b111001111100101101000011, 
24'b000010101101010010111010, 
24'b000000010111101110000001, 
24'b111101010110010000010101, 
24'b000011110001110001110100, 
24'b111100011011001011111101, 
24'b000010001111110110000101, 
24'b111111111000001000011011, 
24'b111101101111111000010111, 
24'b000100001111000111100110, 
24'b111010101110110111111000, 
24'b000101000001001000111010, 
24'b111100101110110110011011, 
24'b000000010001001001110010, 
24'b000011101010110110110101, 
24'b111000001001000111101100, 
24'b001011101111111010101000, 
24'b110001010100000010100011, 
24'b010000010010000000010011, 
24'b101111100111111101010110, 
24'b001111001001000011111100, 
24'b110011000101111100010000, 
24'b001010010100000001111110, 
24'b111000000100000001010011, 
24'b000110010110111010011011, 
24'b111010001010001010001110, 
24'b000110100100110001101000, 
24'b110111101101010001001101, 
24'b001010100101101110000000, 
24'b110011001101010000010110, 
24'b001110010101110011110010, 
24'b110001010101000101111101, 
24'b001101011101000001101011, 
24'b110101010011110110010001, 
24'b000110101100010001000101, 
24'b111110000101101001010011, 
24'b111101000101011001110001, 
24'b000111001011100110000111, 
24'b110101110000010111000100, 
24'b001011110011101110010001, 
24'b110100001110001010110010, 
24'b001010011100111100110110, 
24'b110111110011111100000101, 
24'b000101101110001001011111, 
24'b111100011101110011001010, 
24'b000010010001001101100110, 
24'b111101111001110100001011, 
24'b000011001001000111111100, 
24'b111010111011111101010110, 
24'b000111100001111100110110, 
24'b110110000011001000101100, 
24'b001011110101110010110100, 
24'b110011001111010000010000, 
24'b001100100011101110010001, 
24'b110100110001010001110100, 
24'b001001000110101111001100, 
24'b111001011111001111010010, 
24'b000011111100110010010000, 
24'b111110001101001100101010, 
24'b000000010110110011110010, 
24'b000000010111001100100000, 
24'b111111100100110010101001, 
24'b000000001110001110011011, 
24'b111111111110110000101101, 
24'b000000001110001111101001, 
24'b111110111000110000110111, 
24'b000010101101001101101110, 
24'b111011001001110100100011, 
24'b000111010000001000100110, 
24'b110110100101111010011101, 
24'b001010111010000010101101, 
24'b110100101100111111100100, 
24'b001010011010111111001000, 
24'b110111110011000001001100, 
24'b000100111111111111011110, 
24'b111110110010111111001000, 
24'b111101011110000010101110, 
24'b000101101001111011011011, 
24'b111000010100000110000100, 
24'b001000011000111001001001, 
24'b111000010100000110110010, 
24'b000101110110111010010100, 
24'b111100101001000011101010, 
24'b000000101111111111001011, 
24'b000001011111111101011011, 
24'b111101001000000110010110, 
24'b000011001111110101110010, 
24'b111101011000001101111100, 
24'b000001010011101110101010, 
24'b000000010011010100010000, 
24'b111110010110101001100011, 
24'b000010010101010111110110, 
24'b111101111010100111110011, 
24'b000000111010010111011011, 
24'b000001000000101010100110, 
24'b111100110110010010001000, 
24'b000100111111110010011010, 
24'b111010000111001000000101, 
24'b000101011000111110001000, 
24'b111100101100111011011110, 
24'b111111101111001010100100, 
24'b000100111110110000010111, 
24'b110101111011010011001110, 
24'b001110110001101011001101, 
24'b101101101101010100001011, 
24'b010100000000101110101101, 
24'b101100011111001100100000, 
24'b010000111001111001110001, 
24'b110011100000111111001101, 
24'b000111000100000111101111, 
24'b111110100100110010001111, 
24'b111100101000010010001010, 
24'b000110100110101011101111, 
24'b111000010100010011110111, 
24'b000110100000101111000110, 
24'b111100110001001011110000, 
24'b111110011111111011000101, 
24'b000110111100111101001110, 
24'b110011111010001010011111, 
24'b010000001101101110101010, 
24'b101101011001010110100111, 
24'b010011000011100110010100, 
24'b101110011010011010011001, 
24'b001110100110100111010100, 
24'b110101010001010100111010, 
24'b000110101011110000011010, 
24'b111100110110001001011110, 
24'b000000101111111100101001, 
24'b000000010100111110000010, 
24'b111111111110000101111010, 
24'b111110100111110111111110, 
24'b000011011100001000001000, 
24'b111010011101111001101101, 
24'b000111001110000010111001, 
24'b110111111001000001100100, 
24'b001000000000111001100101, 
24'b111001000000001011000011, 
24'b000101011011110001000111, 
24'b111100010011010001100001, 
24'b000010010010101101001110, 
24'b111110011000010010101010, 
24'b000001111110101110100100, 
24'b111100101001001111011110, 
24'b000101101001110010110100, 
24'b110111100100001011000011, 
24'b001011001111110110101101, 
24'b110010011101001000001010, 
24'b001110111100111000011111, 
24'b110000110111000111010010, 
24'b001110000001111001000000, 
24'b110100001101000110011011, 
24'b001000110001111010110100, 
24'b111010101000000011000111, 
24'b000010000110111111110000, 
24'b000000101010111100110010, 
24'b111101010101000110110111, 
24'b000011110011110101110100, 
24'b111011110100001100101000, 
24'b000100000110110010010011, 
24'b111100001010001101000110, 
24'b000011110011110101010000, 
24'b111011110100000110110111, 
24'b000101001010111110001010, 
24'b111001010101111100010110, 
24'b001000011110001001000000, 
24'b110101101111110010011101, 
24'b001011101011010000110100, 
24'b110011100110101101011111, 
24'b001100001110010010101100, 
24'b110100111100101110011111, 
24'b001001001001001111100000, 
24'b111001010001110010111010, 
24'b000100010010001010110011, 
24'b111101101110110111000011, 
24'b000001001011000111101111, 
24'b111110110101111000110110, 
24'b000010011100000110111010, 
24'b111011001101111001010100, 
24'b000111111101000110001010, 
24'b110100100100111010111111, 
24'b001110101100000011001100, 
24'b101110110010111111010000, 
24'b010010100111111110000011, 
24'b101101010110000100100000, 
24'b010001010101111001101011, 
24'b110001001101000111000000, 
24'b001011011001111001110000, 
24'b111000100000000011111111, 
24'b000011100011111111011110, 
24'b000000000110111100010101, 
24'b111100110100000111111101, 
24'b000101101011110100011000, 
24'b111000011100001110000100, 
24'b001001000000110001001010, 
24'b110101110010001101111011, 
24'b001011010100110100011110, 
24'b110011100100001000010000, 
24'b001101100011111011010010, 
24'b110001011000000001110010, 
24'b001111011010000000000010, 
24'b110000010001111111110010, 
24'b001111011110111110110100, 
24'b110001100010000011111011, 
24'b001100110101111000101010, 
24'b110101010001001010101010, 
24'b001000011100110010111100, 
24'b111001101010001101111001, 
24'b000100110110110011010010, 
24'b111011110100001001100101, 
24'b000100100010111011001001, 
24'b111010001101111111010011, 
24'b000111101111000110001101, 
24'b110110000011110101010100, 
24'b001011111101001101010111, 
24'b110010110111110010010000, 
24'b001101001100001011110010, 
24'b110100001101111000001100, 
24'b001000111111000010100111, 
24'b111011000010000010111001, 
24'b000000010000111000010110, 
24'b000100100101001010110011, 
24'b110111001111110100001101, 
24'b001011101111001010011010, 
24'b110011000001111001000110, 
24'b001100010100000001111011, 
24'b110110001110000011101011, 
24'b000101101011110111001000, 
24'b111111011100001100110110, 
24'b111011000111110001000100, 
24'b001001111110001110110111, 
24'b110001111010110011010010, 
24'b010000110010001000111111, 
24'b101110001110111011101011, 
24'b010001001010111111100111, 
24'b110000111011000100011000, 
24'b001011111110111000111011, 
24'b110111101011001000001010, 
24'b000100100101111000011111, 
24'b111110110111000101100000, 
24'b111110010110111101011101, 
24'b000011101010111111010001, 
24'b111011001100000011110000, 
24'b000101010000111001111110, 
24'b111010110111000111010000, 
24'b000100101000111000101010, 
24'b111100000101000110011010, 
24'b000011001010111011010010, 
24'b111101011110000010101010, 
24'b000010000110111111011001, 
24'b111110000011111110111101, 
24'b000010001001000010000100, 
24'b111101010010111101110001, 
24'b000011110000000001100100, 
24'b111010110000111111111010, 
24'b000111001011111101111101, 
24'b110110100101000100100110, 
24'b001011110011111000101010, 
24'b110001111110001010000101, 
24'b001111110111110011100100, 
24'b101111000111001110001010, 
24'b010000110010110000111011, 
24'b110000101000001110111111, 
24'b001100100011110010001101, 
24'b110111100101001011100010, 
24'b000011010001110111101000, 
24'b000010100010000100101001, 
24'b110111100111111111001011, 
24'b001101110000111101011011, 
24'b101101111011000101000001, 
24'b010100111101111001111110, 
24'b101001111001000101010111, 
24'b010101100101111101000010, 
24'b101100100010111111000110, 
24'b010000001010000101101111, 
24'b110011111010110101001011, 
24'b000111101111001111011010, 
24'b111100011101101101010100, 
24'b111111111010010100001011, 
24'b000011000011101100011001, 
24'b111010110001010001001000, 
24'b000110101110110010110001, 
24'b111000010111001000101111, 
24'b001000001101111011011110, 
24'b110111011010000001100101, 
24'b001000111010111111011011, 
24'b110110110011000001111101, 
24'b001001011110111010011111, 
24'b110110011011001010110101, 
24'b001001100100101111000011, 
24'b110110110000010110110000, 
24'b001000101101100100111000, 
24'b111000000000011101000110, 
24'b000111010000100011110101, 
24'b111001011010011000010000, 
24'b000110001111101110001001, 
24'b111001110000001001111010, 
24'b000110101100111110011001, 
24'b111000100100111010010001, 
24'b001000011000001011000001, 
24'b110110110111110010100001, 
24'b001001100001001100110101, 
24'b110110110111110110101100, 
24'b000111110111000011110000, 
24'b111010011011000010110110, 
24'b000010010111110110110011, 
24'b000001100010001110010000, 
24'b111010001101101110110010, 
24'b001001111110010001101111, 
24'b110010011000110000000110, 
24'b010000011001001100010100, 
24'b101110000000111000001100, 
24'b010010011000000011010111, 
24'b101110011111000000001000, 
24'b001111101011111101111111, 
24'b110010110111000010000100, 
24'b001010010000111111100010, 
24'b111000101010111101100111, 
24'b000100110001000101101100, 
24'b111101010011110111010100, 
24'b000001001110001010110000, 
24'b111111101010110100100001, 
24'b111111111101001010110011, 
24'b000000000101110111000011, 
24'b000000000110000110011110, 
24'b111111101100111100000001, 
24'b000000011111000010001001, 
24'b111111011111111110101001, 
24'b000000011110000001110010, 
24'b111111101111111100101110, 
24'b000000000010000101011011, 
24'b000000001110111000011010, 
24'b111111100110001001001001, 
24'b000000100100110110011100, 
24'b111111010110001000100100, 
24'b000000101100111001110011, 
24'b111111010110000010110101, 
24'b000000100111000000111011, 
24'b111111011110111011101011, 
24'b000000011110000110101011, 
24'b111111100100111000101011, 
24'b000000011100000110001010, 
24'b111111011110111100110001, 
24'b000000101111111111000010, 
24'b111111000000000101101111, 
24'b000001010111110101110010, 
24'b111110010001001101101010, 
24'b000010000011110000100101, 
24'b111101110111001111010010, 
24'b000001111011110010101001, 
24'b111110110100001010000010, 
24'b111111110111111010000011, 
24'b000010000110000001111011, 
24'b111011011000000001011010, 
24'b000111100100111100011101, 
24'b110101011000000100011000, 
24'b001101100010111011111111, 
24'b110000001001000010111100, 
24'b010001010011111110001101, 
24'b101110011010000001001110, 
24'b010000101000111110001101, 
24'b110001100011000011110011, 
24'b001011010010111000110011, 
24'b111000011101001011101000, 
24'b000011101011101111100010, 
24'b111111110111010100111010, 
24'b111101010110100111111010, 
24'b000100011010011001011010, 
24'b111011000001100111100010, 
24'b000100100011010101010010, 
24'b111100101001101111110110, 
24'b000001110010001001110010, 
24'b111111101101111100111111, 
24'b111111010011111100101110, 
24'b000000111010001000010001, 
24'b111111110000110100100110, 
24'b111110101111001100011010, 
24'b000011010100110100100111, 
24'b111010011101001000101111, 
24'b000111100000111010111110, 
24'b110111001111000000111101, 
24'b001001000000000010110101, 
24'b110111111001111010001101, 
24'b000110000100000111100111, 
24'b111100111101110111110000, 
24'b111111011000000111110101, 
24'b000100100011111001010100, 
24'b110111101000000101001101, 
24'b001011101111111100001111, 
24'b110001100101000010101101, 
24'b010000010110111101110100, 
24'b101110011101000010001111, 
24'b010010000000111101001110, 
24'b101110001001000011100101, 
24'b010001001011111011100101, 
24'b101111111110000101000100, 
24'b001110011000111010101101, 
24'b110011110010000101000111, 
24'b001001011111111011100011, 
24'b111001110001000011011100, 
24'b000010100101111101110010, 
24'b000001010011000000111011, 
24'b111010111111000000001100, 
24'b001000001101111110111011, 
24'b110101100010000001100111, 
24'b001011011111111110001011, 
24'b110100111100000001101111, 
24'b001001001110111110100100, 
24'b111001110110000001000110, 
24'b000010010111111111010001, 
24'b000001100101000000100001, 
24'b111010111111111111100001, 
24'b000111010110000000101100, 
24'b110111111001111110111011, 
24'b000111000111000001100111, 
24'b111011100011111101110010, 
24'b000000011100000010110000, 
24'b000100010000111100111100, 
24'b110111000011000011000001, 
24'b001100111011111101011110, 
24'b110000011111000001100001, 
24'b010000011001000000000011, 
24'b110000100110111110000000, 
24'b001100110000000100001101, 
24'b110111001011111001101000, 
24'b000100010000001000010000, 
24'b000000010100110110100100, 
24'b111011101011001001101111, 
24'b000111011000110111000101, 
24'b110110110011000110111111, 
24'b001001110111111100000001, 
24'b110110011110000000010011, 
24'b001000100100000011101110, 
24'b111000101010111000011100, 
24'b000110001100001010101101, 
24'b111010110000110011010011, 
24'b000100101000001101001110, 
24'b111011111001110011110100, 
24'b000011100011001001110000, 
24'b111101011000111001110001, 
24'b000001001001000010000111, 
24'b0_00001000101000001111110, 
24'b001111010001000100001011, 
24'b110001000010111100010100, 
24'b001110011101000011000010, 
24'b110010010001111101110001, 
24'b001100110110000001010010, 
24'b110100001101111111110001, 
24'b001010101000111111000100, 
24'b110110100111000010001100, 
24'b001000000111111100100010, 
24'b111001001011000100110011, 
24'b000101100011111001111000, 
24'b111011101001000111011000, 
24'b000011010000110111011010, 
24'b111101101101001001101110, 
24'b000001011110110101010010, 
24'b111111001000001011100101, 
24'b000000011101110011101110, 
24'b111111101111001100110010, 
24'b000000010011110010111011, 
24'b111111011011001101001100, 
24'b000001000111110010111011, 
24'b111110001010001100101111, 
24'b000010110011110011110101, 
24'b111100000010001011011010, 
24'b000101010100110101100011, 
24'b111001001100001001010100, 
24'b001000011100111000000001, 
24'b110101110110000110100010, 
24'b001011111010111011000011, 
24'b110010010100000011010010, 
24'b001111011011111110011101, 
24'b101110110111111111110010, 
24'b010010101110000001111110, 
24'b101011110011111100010011, 
24'b010101011111000101011000, 
24'b101001011100111001000010, 
24'b010111011100001000011100, 
24'b100111111100110110001111, 
24'b011000011011001010111100, 
24'b100111011111110100000100, 
24'b011000010100001100101111, 
24'b101000001001110010101001, 
24'b010111001000001101110000, 
24'b101001110110110010000011, 
24'b010100111010001101111011, 
24'b101100100001110010010011, 
24'b010001110101001101010110, 
24'b101111111110110011001110, 
24'b001110000110001100000100, 
24'b110011111011110100110100, 
24'b001010000001001010001111, 
24'b111000000100110110110101, 
24'b000101111010001000000011, 
24'b111100000110111001000110, 
24'b000010000000000101101101, 
24'b111111101111111011011110, 
24'b111110101010000011011010, 
24'b000010110010111101101101, 
24'b111100000010000001010010, 
24'b000100111101111111101010, 
24'b111010010100111111100000, 
24'b000110001100000001001111, 
24'b111001100100111110001001, 
24'b000110011100000010010111, 
24'b111001110010111101010001, 
24'b000101110100000011000000, 
24'b111010110100111100110111, 
24'b000100011000000011001100, 
24'b111100100011111100110111, 
24'b000010011010000011000001, 
24'b111110101111111101001010, 
24'b000000000110000010100101, 
24'b000001001000111101101011, 
24'b111101101101000010000011, 
24'b000011011101111110010000, 
24'b111011100001000001011110, 
24'b000101011100111110110001, 
24'b111001110000000001000011, 
24'b000110111011111111000110, 
24'b111000100101000000110101, 
24'b000111101110111111001011, 
24'b111000001001000000111010, 
24'b000111110001111110111100, 
24'b111000100000000001010011, 
24'b000111000101111110011001, 
24'b111001100101000010000000, 
24'b000101101010111101100100, 
24'b111011010000000010111011, 
24'b000011101101111100100011, 
24'b111101011011000011111111, 
24'b000001011001111011011110, 
24'b111111110110000101000101, 
24'b111110111011111010011000, 
24'b000010010101000110000101, 
24'b111100011111111001011111, 
24'b000100101001000110110101, 
24'b111010010100111000111010, 
24'b000110100111000111001110, 
24'b111000100101111000101111, 
24'b001000000100000111001010, 
24'b110111011010111001000100, 
24'b001000111101000110100101, 
24'b110110110101111001111011, 
24'b001001001111000101011100, 
24'b110110110110111011010101, 
24'b001000111101000011110010, 
24'b110111011001111101010001, 
24'b001000001011000001101000, 
24'b111000010110111111100111, 
24'b000111000110111111000100, 
24'b111001100010000010010110, 
24'b000101110101111100001110, 
24'b111010110001000101010000, 
24'b000100101000111001001111, 
24'b111011111011001000010010, 
24'b000011100110110110001111, 
24'b111100110011001011010001, 
24'b000010111011110011010100, 
24'b111101010001001110000101, 
24'b000010101011110000101000, 
24'b111101010001010000100110, 
24'b000010111001101110010000, 
24'b111100110100010010110010, 
24'b000011100101101100010001, 
24'b111011111100010100100110, 
24'b000100100110101010101101, 
24'b111010110001010101111101, 
24'b000101111000101001100010, 
24'b111001011101010110111001, 
24'b000111001110101000110010, 
24'b111000001000010111011100, 
24'b001000011101101000011011, 
24'b110111000011010111100111, 
24'b001001011000101000011011, 
24'b110110010110010111011110, 
24'b001001110010101000101011, 
24'b110110001110010111000100, 
24'b001001100111101001001110, 
24'b110110101110010110011010, 
24'b001000110000101001111111, 
24'b110111111100010101100011, 
24'b000111001101101010111101, 
24'b111001110100010100011111, 
24'b000101000001101100001000, 
24'b111100010011010011001101, 
24'b000010010011101101100010, 
24'b111111001101010001101100, 
24'b111111001111101111001011, 
24'b000010010110001111111010, 
24'b111100000011110001000101, 
24'b000101100001001101110110, 
24'b111001000000110011010010, 
24'b001000011011001011100000, 
24'b110110010010110101110010, 
24'b001010111001001000110101, 
24'b110100000111111000101000, 
24'b001100101110000101111000, 
24'b110010101010111011101101, 
24'b001101110000000010101001, 
24'b110010000101111111000011, 
24'b001101111001111111001111, 
24'b110010011000000010100001, 
24'b001101001001111011101110, 
24'b110011100011000110000010, 
24'b001011100100111000001111, 
24'b110101100000001001011101, 
24'b001001001111110100111011, 
24'b111000001000001100101000, 
24'b000110011010110001111100, 
24'b111011001010001111011010, 
24'b000011001101101111011000, 
24'b111110011011010001101001, 
24'b111111111100101101100001, 
24'b000001101010010011001010, 
24'b111100110011101100010110, 
24'b000100101001010011111011, 
24'b111010000001101100000011, 
24'b000111001101010011110001, 
24'b110111101110101100101010, 
24'b001001001101010010101110, 
24'b110110000100101110001000, 
24'b001010100001010000110100, 
24'b110101000100110000011100, 
24'b001011001010001110000110, 
24'b110100110001110011100000, 
24'b001011001010001010101110, 
24'b110101000100110111001011, 
24'b001010100100000110110101, 
24'b110101111001111011001111, 
24'b001001100011000010101011, 
24'b110111000100111111011101, 
24'b001000010001111110011100, 
24'b111000011011000011101000, 
24'b000110111000111010011010, 
24'b111001110100000111011110, 
24'b000101100010110110110011, 
24'b111011000011001010110001, 
24'b000100011010110011110110, 
24'b111100000101001101010101, 
24'b000011100010110001101110, 
24'b111100110001001110111110, 
24'b000011000010110000100110, 
24'b111101000110001111100110, 
24'b000010110111110000011111, 
24'b111101000110001111001001, 
24'b000011000001110001011110, 
24'b111100110100001101101011, 
24'b000011011001110011011100, 
24'b111100011000001011001110, 
24'b000011110111110110010101, 
24'b111011111010000111111110, 
24'b000100010011111001111011, 
24'b111011100010000100000100, 
24'b000100100100111110000011, 
24'b111011011010111111110010, 
24'b000100100100000010011010, 
24'b111011100101111011011010, 
24'b000100001011000110110000, 
24'b111100001010110111001100, 
24'b000011010111001010110001, 
24'b111101001101110011011011, 
24'b000010001000001110001101, 
24'b111110101010110000010111, 
24'b000000011111010000110111, 
24'b000000011101101110001101, 
24'b111110100011010010011111, 
24'b000010011110101101001000, 
24'b111100011110010010111111, 
24'b000100100110101101001110, 
24'b111010010111010010010010, 
24'b000110101001101110100010, 
24'b111000011101010000011000, 
24'b001000011001110001000001, 
24'b110110110111001101010110, 
24'b001001101111110100100011, 
24'b110101110011001001010101, 
24'b001010100001111001000000, 
24'b110101010110000100100010, 
24'b001010101000111110000110, 
24'b110101100111111111001101, 
24'b001010000000000011100110, 
24'b110110100101111001100110, 
24'b001000101001001001001110, 
24'b111000010100110100000011, 
24'b000110100101001110101000, 
24'b111010101100101110110100, 
24'b000011111101010011100100, 
24'b111101100100101010001111, 
24'b000000110101010111101111, 
24'b000000110101100110100010, 
24'b111101011110011010111011, 
24'b000100010010100011111010, 
24'b111001111110011100111110, 
24'b000111101110100010100000, 
24'b110110100111011101101110, 
24'b001011000000100010011001, 
24'b110011100000011101001010, 
24'b001101111001100011100111, 
24'b110000110100011011010100, 
24'b010000010100100110000011, 
24'b101110101100011000010010, 
24'b010010001001101001101001, 
24'b101101001011010100001110, 
24'b010011010110101110001000, 
24'b101100010011001111010110, 
24'b010011111001110011010101, 
24'b101100000100001001111001, 
24'b010011110101111000111101, 
24'b101100011001000100001011, 
24'b010011010001111110101101, 
24'b101101001110111110011100, 
24'b010010010001000100010100, 
24'b101110010111111001000001, 
24'b010000111110001001100010, 
24'b101111110000110100000111, 
24'b001111100010001110000100, 
24'b110001001110101111111111, 
24'b001110000010010001110000, 
24'b110010101010101100110011, 
24'b001100101011010100011011, 
24'b110011111111101010101011, 
24'b001011011101010101111110, 
24'b110101000100101001101010, 
24'b001010100001010110011100, 
24'b110101111000101001101110, 
24'b001001110110010101110101, 
24'b110110011001101010110110, 
24'b001001011101010100001111, 
24'b110110100111101100110111, 
24'b001001010110010001110101, 
24'b110110100111101111101001, 
24'b001001011101001110110011, 
24'b110110011101110010111011, 
24'b001001101011001011010101, 
24'b110110001010110110100000, 
24'b001001111111000111101100, 
24'b110101111001111010001000, 
24'b001010001110000100000110, 
24'b110101101011111101100111, 
24'b001010011001000000110010, 
24'b110101100111000000101110, 
24'b001010010110111101111100, 
24'b110101110001000011010000, 
24'b001010000110111011101110, 
24'b110110001010000101001000, 
24'b001001100011111010001111, 
24'b110110110101000110001101, 
24'b001000110000111001100100, 
24'b110111110010000110011111, 
24'b000111101010111001101011, 
24'b111000111110000101111111, 
24'b000110010111111010100001, 
24'b111010011000000100110011, 
24'b000100110111111100000001, 
24'b111011111100000011000010, 
24'b000011010000111110000010, 
24'b111101100110000000110101, 
24'b000001100101000000011000, 
24'b111111010001111110011001, 
24'b111111111100000010110110, 
24'b000000111000111011111011, 
24'b111110011000000101010001, 
24'b000010010111111001100110, 
24'b111100111110000111011011, 
24'b000011101100110111101000, 
24'b111011110000001001001011, 
24'b000100110001110110001011, 
24'b111010110000001010010101, 
24'b000101101010110101010110, 
24'b111010000001001010110011, 
24'b000110010011110101001111, 
24'b111001011111001010100001, 
24'b000110101100110101111000, 
24'b111001001100001001100011, 
24'b000110111010110111001111, 
24'b111001000010000111110111, 
24'b000110111111111001001111, 
24'b111001000010000101100101, 
24'b000110111110111011110000, 
24'b111001000100000010110111, 
24'b000110111100111110101001, 
24'b111001000100111111111000, 
24'b000110111110000001101010, 
24'b111000111110111100110101, 
24'b000111000111000100101001, 
24'b111000110000111001111110, 
24'b000111011011000111010111, 
24'b111000010110110111011101, 
24'b000111111110001001100111, 
24'b110111101100110101100000, 
24'b001000110000001011001100, 
24'b110110110010110100010010, 
24'b001001110001001100000011, 
24'b110101101010110011111001, 
24'b001011000001001011111110, 
24'b110100010010110100011001, 
24'b001100011101001011000011, 
24'b110010110001110101110001, 
24'b001110000001001001001111, 
24'b110001001100110111111101, 
24'b001111101000000110101100, 
24'b101111100110111010110111, 
24'b010001001010000011100000, 
24'b101110001000111110010001, 
24'b010010100011111111111001, 
24'b101100110111000010000000, 
24'b010011101010111100000110, 
24'b101011111100000101110011, 
24'b010100011001111000010111, 
24'b101011011001001001011011, 
24'b010100101101110100111100, 
24'b101011010110001100100111, 
24'b010100011111110010000010, 
24'b101011110011001111001100, 
24'b010011110001101111110110, 
24'b101100110011010000111100, 
24'b010010100000101110100000, 
24'b101110010011010001110101, 
24'b010000110001101110000111, 
24'b110000010001010001110000, 
24'b001110100110101110101000, 
24'b110010100110010000110000, 
24'b001100001010110000000101, 
24'b110101001011001110111011, 
24'b001001011111110010010000, 
24'b110111111001001100011010, 
24'b000110110011110101000001, 
24'b111010100010001001011101, 
24'b000100001100111000001000, 
24'b111101000011000110010001, 
24'b000001110101111011010100, 
24'b111111001110000011001001, 
24'b111111110101111110010110, 
24'b000001000000000000010010, 
24'b111110010100000000111101, 
24'b000010010010111101111101, 
24'b111101010001000010111110, 
24'b000011000010111100010100, 
24'b111100110011000100001011, 
24'b000011001111111011100011, 
24'b111100110101000100100010, 
24'b000010111101111011101001, 
24'b111101010111000011111110, 
24'b000010010000111100100111, 
24'b111110001101000010100101, 
24'b000001010010111110011000, 
24'b111111010010000000100000, 
24'b000000001000000000110010, 
24'b000000011111111101111000, 
24'b111110111100000011100100, 
24'b000001100101111010111110, 
24'b111101111011000110100010, 
24'b000010100000111000000001, 
24'b111101001010001001011001, 
24'b000011000101110101010010, 
24'b111100110011001011111100, 
24'b000011001111110011000010, 
24'b111100111000001101110111, 
24'b000010111010110001011100, 
24'b111101011100001111000101, 
24'b000010000101110000101010, 
24'b111110100000001111011010, 
24'b000000110101110000110000, 
24'b111111111101001110110111, 
24'b111111001011110001101110, 
24'b000001110000001101011110, 
24'b111101010000110011100000, 
24'b000011110000001011011000, 
24'b111011001101110101111100, 
24'b000101110100001000101101, 
24'b111001001101111000110000, 
24'b000111110000000101110000, 
24'b110111010111111011110001, 
24'b001001011100000010110000, 
24'b110101111000111110101011, 
24'b001010101110111111111111, 
24'b110100110100000001001111, 
24'b001011100001111101101011, 
24'b110100010100000011001101, 
24'b001011110001111100000110, 
24'b110100010110000100011010, 
24'b001011011010111011010100, 
24'b110100111101000100101111, 
24'b001010100011111011011110, 
24'b110110000101000100001000, 
24'b001001001011111100100000, 
24'b110111101001000010101001, 
24'b000111011110111110011000, 
24'b111001011111000000011101, 
24'b000101100010000000111000, 
24'b111011011111111101101101, 
24'b000011100001000011110010, 
24'b111101011110111010101100, 
24'b000001100111000110110111, 
24'b111111010010110111101001, 
24'b111111111010001001110010, 
24'b000000110011110100111001, 
24'b111110100110001100010011, 
24'b000001111010110010101101, 
24'b111101101110001110001000, 
24'b000010100010110001010001, 
24'b111101010111001111000110, 
24'b000010101001110000110011, 
24'b111101011111001111000100, 
24'b000010010000110001010111, 
24'b111110001001001101111101, 
24'b000001011010110010111111, 
24'b111111001010001011110110, 
24'b000000001110110101100011, 
24'b000000100000001000110110, 
24'b111110101111111000111011, 
24'b000010000001000101001001, 
24'b111101001100111100111001, 
24'b000011101000000001000000, 
24'b111011101000000001001011, 
24'b000101000110111100101100, 
24'b111010001101000101011110, 
24'b000110011011111000011110, 
24'b111001000010001001011111, 
24'b000111011011110100101101, 
24'b111000001111001100111101, 
24'b001000000010110001100110, 
24'b110111110101001111101010, 
24'b001000001110101111010110, 
24'b110111110110010001011100, 
24'b001000000000101110000010, 
24'b111000010000010010001110, 
24'b000111011000101101110010, 
24'b111001000101010001111111, 
24'b000110011000101110011110, 
24'b111010001101010000110100, 
24'b000101001000110000000101, 
24'b111011100110001110110111, 
24'b000011101000110010011000, 
24'b111101001001001100010010, 
24'b000010000100110101001010, 
24'b111110101111001001010101, 
24'b000000011100111000001110, 
24'b000000010110000110001110, 
24'b111110111001111011010001, 
24'b000001110111000011010000, 
24'b111101011100111110000111, 
24'b000011001101000000100101, 
24'b111100001010000000100100, 
24'b000100011010111110011001, 
24'b111011000110000010011101, 
24'b000101010111111100110100, 
24'b111010010000000011101111, 
24'b000110000110111011111000, 
24'b111001100110000100010111, 
24'b000110100111111011100011, 
24'b111001001100000100010111, 
24'b000110111100111011110101, 
24'b111000111110000011110110, 
24'b000111000101111100100101, 
24'b111000111011000010111010, 
24'b000111000010111101101010, 
24'b111001000100000001101111, 
24'b000110110101111110111011, 
24'b111001010011000000011100, 
24'b000110100001000000001100, 
24'b111001101101111111001101, 
24'b000110000011000001011001, 
24'b111010001100111110000111, 
24'b000101100010000010010110, 
24'b111010110001111101010010, 
24'b000100111000000011000000, 
24'b111011011100111100110011, 
24'b000100001101000011010110, 
24'b111100001001111100100111, 
24'b000011100000000011010111, 
24'b111100110111111100110000, 
24'b000010110011000011001000, 
24'b111101100011111101000111, 
24'b000010001000000010101000, 
24'b111110001011111101101011, 
24'b000001100101000010000000, 
24'b111110101010111110010101, 
24'b000001001011000001010101, 
24'b111110111111111111000000, 
24'b000000111101000000101100, 
24'b111111000011111111100110, 
24'b000001000000000000001000, 
24'b111110111000000000000110, 
24'b000001010110111111101110, 
24'b111110011000000000011100, 
24'b000010000000111111011100, 
24'b111101100100000000101010, 
24'b000010111101111111010100, 
24'b111100011110000000101111, 
24'b000100001100111111010001, 
24'b111011001000000000101111, 
24'b000101101010111111010001, 
24'b111001100100000000101111, 
24'b000111010011111111010001, 
24'b110111110111000000110010, 
24'b001000111111111111001011, 
24'b110110001100000000111001, 
24'b001010101000111111000000, 
24'b110100100111000001001010, 
24'b001100000111111110101011, 
24'b110011010001000001100011, 
24'b001101010011111110001110, 
24'b110010010000000010000100, 
24'b001110000110111101100111, 
24'b110001101010000010101110, 
24'b001110011101111100111110, 
24'b110001100101000011011001, 
24'b001110010010111100010001, 
24'b110010000010000100000100, 
24'b001101100010111011101010, 
24'b110011000000000100100110, 
24'b001100010101111011001010, 
24'b110100011111000100111111, 
24'b001010100111111010111000, 
24'b110110011001000101001001, 
24'b001000100010111010111000, 
24'b111000100111000101000001, 
24'b000110001110111011001010, 
24'b111010111111000100100110, 
24'b000011110100111011101101, 
24'b111101011001000011111011, 
24'b000001011100111100100000, 
24'b111111101101000011000010, 
24'b111111001111111101011110, 
24'b000001101110000010000001, 
24'b111101011001111110100010, 
24'b000011011001000000111110, 
24'b111011111100111111100001, 
24'b000100100110000000000001, 
24'b111011000001000000011001, 
24'b000101010001111111010010, 
24'b111010100101000000111110, 
24'b000101011100111110111000, 
24'b111010101010000001001110, 
24'b000101001000111110110101, 
24'b111011001111000001000001, 
24'b000100010110111111010001, 
24'b111100001101000000011001, 
24'b000011001100000000000110, 
24'b111101011111111111010100, 
24'b000001110011000001010111, 
24'b111110111111111101111001, 
24'b000000001111000010111101, 
24'b000000100100111100001100, 
24'b111110101001000100101111, 
24'b000010001011111010010110, 
24'b111101000010000110100101, 
24'b000011101111111000100001, 
24'b111011100010001000010111, 
24'b000101001101110110110110, 
24'b111010001000001001111000, 
24'b000110100011110101011111, 
24'b111000110100001011000100, 
24'b000111110100110100100010, 
24'b110111100101001011110001, 
24'b001001000010110100000100, 
24'b110110011000001011111101, 
24'b001010001111110100001010, 
24'b110101001000001011100101, 
24'b001011100001110100110010, 
24'b110011110010001010101111, 
24'b001100111101110101110110, 
24'b110010010011001001011111, 
24'b001110100001110111010010, 
24'b110000100110000111111011, 
24'b010000010100111000111011, 
24'b101110101111000110001101, 
24'b010010010001111010101010, 
24'b101100101110000100011111, 
24'b010100010110111100010100, 
24'b101010100110000010111101, 
24'b010110011101111101101101, 
24'b101000011111000001101110, 
24'b011000100001111110110010, 
24'b100110100010000000110110, 
24'b011010010110111111011001, 
24'b100100111000000000011101, 
24'b011011110100111111100111, 
24'b100011101000000000011111, 
24'b011100110001111111010101, 
24'b100010111110000000111101, 
24'b011101000111111110101101, 
24'b100010111110000001101111, 
24'b011100101110111101110001, 
24'b100011110000000010110000, 
24'b011011100110111100101101, 
24'b100101010001000011110110, 
24'b011001101011111011101000, 
24'b100111100011000100111000, 
24'b010111000100111010101010, 
24'b101010011101000101101111, 
24'b010011111000111001111101, 
24'b101101110111000110010011, 
24'b010000010001111001100100, 
24'b110001100110000110011111, 
24'b001100011110111001100100, 
24'b110101011010000110010011, 
24'b001000101101111001111010, 
24'b111001001000000101110011, 
24'b000101001010111010100101, 
24'b111100011100000101000001, 
24'b000010000100111011011011, 
24'b111111001111000100000101, 
24'b111111100111111100011000, 
24'b000001010110000011001001, 
24'b111101111001111101010001, 
24'b000010101000000010010111, 
24'b111101000010111101111101, 
24'b000011000101000001110101, 
24'b111100111110111110010010, 
24'b000010110000000001101100, 
24'b111101101011111110001110, 
24'b000001101111000010000001, 
24'b111111000000111101101001, 
24'b000000001011000010110100, 
24'b000000101111111100100111, 
24'b111110010001000100000100, 
24'b000010101111111011001100, 
24'b111100010001000101101010, 
24'b000100101101111001011110, 
24'b111010011000000111011110, 
24'b000110011110110111101000, 
24'b111000110100001001010001, 
24'b000111110000110101111000, 
24'b110111110101001010111010, 
24'b001000011101110100011011, 
24'b110111011101001100001011, 
24'b001000011101110011011011, 
24'b110111110011001100110110, 
24'b000111101110110011000110, 
24'b111000111010001100110011, 
24'b000110010011110011100000, 
24'b111010101100001011111110, 
24'b000100001111110100110001, 
24'b111100111111001010010100, 
24'b000001101110110110110101, 
24'b111111101011000111111001, 
24'b111110111001111001100100, 
24'b000010100010000100110110, 
24'b111100000010111100111000, 
24'b000101010111000001010101, 
24'b111001010011000000100001, 
24'b000111111100111101100111, 
24'b110110111010000100001111, 
24'b001010000110111001111110, 
24'b110101000011000111110000, 
24'b001011101011110110101010, 
24'b110011110001001010110011, 
24'b001100100111110011111011, 
24'b110011001011001101001011, 
24'b001100110110110001111110, 
24'b110011010001001110101011, 
24'b001100011101110000111110, 
24'b110011111101001111001011, 
24'b001011100000110000111111, 
24'b110101001010001110101001, 
24'b001010000111110001111111, 
24'b110110101100001101001011, 
24'b001000011111110011111001, 
24'b111000011001001010110110, 
24'b000110110000110110100100, 
24'b111010000110000111111001, 
24'b000101001000111001101101, 
24'b111011101000000100100101, 
24'b000011101111111101001010, 
24'b111100110101000001001010, 
24'b000010101111000000100001, 
24'b111101100111111101111000, 
24'b000010001001000011101001, 
24'b111101111101111010111111, 
24'b000010000100000110001110, 
24'b111101110100111000101111, 
24'b000010011010001000001010, 
24'b111101010001110111001100, 
24'b000011001000001001010001, 
24'b111100011010110110011110, 
24'b000100000110001001100110, 
24'b111011010101110110100011, 
24'b000101001111001001001010, 
24'b111010001101110111010101, 
24'b000110010101001000000110, 
24'b111001001011111000101000, 
24'b000111010011000110100110, 
24'b111000010110111010010000, 
24'b000111111110000100110111, 
24'b110111110101111100000010, 
24'b001000010010000011001000, 
24'b110111101100111101101011, 
24'b001000001101000001100100, 
24'b111000000000111111000011, 
24'b000111101110000000011100, 
24'b111000101001111111111101, 
24'b000110111000111111110010, 
24'b111001101011000000010101, 
24'b000101101111111111101110, 
24'b111010111011000000000110, 
24'b000100011000000000001110, 
24'b111100010100111111010110, 
24'b000011000000000001001100, 
24'b111101101101111110001011, 
24'b000001101000000010100000, 
24'b111111000000111100110001, 
24'b000000011100000011111110, 
24'b000000000110111011010011, 
24'b111111011111000101011000, 
24'b000000111001111001111111, 
24'b111110110101000110100001, 
24'b000001011001111001000100, 
24'b111110011111000111001110, 
24'b000001100100111000101001, 
24'b111110011111000111010100, 
24'b000001011100111000111001, 
24'b111110101110000110101110, 
24'b000001000101111001110100, 
24'b111111001010000101011100, 
24'b000000100101111011011100, 
24'b111111101011000011100010, 
24'b000000000100111101100111, 
24'b000000001100000001000111, 
24'b111111100110000000001111, 
24'b000000100111111110010110, 
24'b111111001111000011000100, 
24'b000000110110111011100010, 
24'b111111000111000101110111, 
24'b000000111001111000110110, 
24'b111111001011001000011000, 
24'b000000101110110110100011, 
24'b111111011101001010011001, 
24'b000000011000110100111000, 
24'b111111110110001011101110, 
24'b111111111010110011111011, 
24'b000000010011001100001111, 
24'b111111011101110011110101, 
24'b000000101111001011111001, 
24'b111111001000110100100111, 
24'b000000111101001010101110, 
24'b111111000010110110001011, 
24'b000000111010001000110010, 
24'b111111010010111000011010, 
24'b000000011100000110010100, 
24'b000000000000111011000011, 
24'b111111011101000011100001, 
24'b000001001110111101111100, 
24'b111101111101000000101000, 
24'b000011000000000000110001, 
24'b111011111100111101111100, 
24'b000101010000000011010000, 
24'b111001011101111011101101, 
24'b000111111011000101001101, 
24'b110110101000111010000101, 
24'b001010111000000110011011, 
24'b110011100111111001010010, 
24'b001101111010000110110101, 
24'b110000100110111001010100, 
24'b010000110101000110010101, 
24'b101101110011111010001101, 
24'b010011011101000101000010, 
24'b101011011010111011111000, 
24'b010101100100000011000010, 
24'b101001101011111110001011, 
24'b010110111100000000100000, 
24'b101000101101000000111000, 
24'b010111011100111101101101, 
24'b101000101010000011101111, 
24'b010111000000111010110111, 
24'b101001100110000110011111, 
24'b010101100111111000010000, 
24'b101011011101001000111011, 
24'b010011010001110110000100, 
24'b101110001111001010110010, 
24'b010000000110110100100011, 
24'b110001101110001011111100, 
24'b001100010011110011110010, 
24'b110101110010001100010010, 
24'b001000000100110011110110, 
24'b111010001011001011110011, 
24'b000011101000110100101111, 
24'b111110100110001010100011, 
24'b111111010001110110011000, 
24'b000010110010001000100111, 
24'b111011010001111000100100, 
24'b000110100011000110001010, 
24'b110111110110111011001100, 
24'b001001100111000011011011, 
24'b110101001011111101111111, 
24'b001011110110000000100101, 
24'b110011011011000000110011, 
24'b001101000111111101110111, 
24'b110010101001000011011010, 
24'b001101011001111011011010, 
24'b110010110101000101101010, 
24'b001100101100111001011001, 
24'b110011111111000111011100, 
24'b001011001010110111110111, 
24'b110101111001001000101011, 
24'b001000111000110110111001, 
24'b111000011110001001011001, 
24'b000110000101110110011101, 
24'b111011011100001001100110, 
24'b000010111110110110011101, 
24'b111110100111001001011001, 
24'b111111110100110110110110, 
24'b000001101111001000111001, 
24'b111100110011110111011100, 
24'b000100100110001000001101, 
24'b111010001000111000001011, 
24'b000111000010000111011110, 
24'b111000000000111000111010, 
24'b001000110110000110110000, 
24'b110110011110111001100101, 
24'b001010000001000110001000, 
24'b110101101010111010001001, 
24'b001010011111000101101000, 
24'b110101100100111010100110, 
24'b001010010001000101001101, 
24'b110110000101111010111110, 
24'b001001011100000100110111, 
24'b110111001011111011010101, 
24'b001000001001000100011011, 
24'b111000101011111011110101, 
24'b000110011111000011110110, 
24'b111010011101111100100011, 
24'b000100101001000010111101, 
24'b111100010001111101100111, 
24'b000010110100000001101011, 
24'b111110000100111111001000, 
24'b000001001010111111111100, 
24'b111111100110000001001000, 
24'b111111110001111101101011, 
24'b000000110011000011101001, 
24'b111110110001111010111010, 
24'b000001100011000110101001, 
24'b111110010001110111101100, 
24'b000001110101001010000100, 
24'b111110001110110100000111, 
24'b000001101000001101110000, 
24'b111110101010110000010111, 
24'b000000111110010001100010, 
24'b111111011111101100100111, 
24'b111111111101010101001101, 
24'b000000101010101001000100, 
24'b111110101011011000100100, 
24'b000010000011100101111100, 
24'b111101010001011011011010, 
24'b000011011110100011011011, 
24'b111011110100011101100100, 
24'b000100111000100001101011, 
24'b111010011111011110111000, 
24'b000110001000100000110011, 
24'b111001010110011111010010, 
24'b000111000110100000111001, 
24'b111000100010011110101101, 
24'b000111110000100001111100, 
24'b111000000100011101001110, 
24'b001000000011100011110111, 
24'b110111111101011010111000, 
24'b000111111100100110100101, 
24'b111000001111010111110110, 
24'b000111100010101001111001, 
24'b111000110011010100010001, 
24'b000110110101101101101011, 
24'b111001100110010000010101, 
24'b000101111110110001101100, 
24'b111010100001001100010010, 
24'b000101000001110101110001, 
24'b111011011110001000010000, 
24'b000100000110111001101101, 
24'b111100010100000100011011, 
24'b000011010110111101011000, 
24'b111100111110000000111010, 
24'b000010110110000000101011, 
24'b111101010010111101110111, 
24'b000010101001000011100001, 
24'b111101010100111011001111, 
24'b000010110110000101111000, 
24'b111100111011111001001001, 
24'b000011011011000111110000, 
24'b111100001010110111011110, 
24'b000100010110001001001101, 
24'b111011000110110110001111, 
24'b000101100011001010001111, 
24'b111001110000110101011000, 
24'b000110111110001010111101, 
24'b111000010011110100110010, 
24'b001000011101001011011010, 
24'b110110110101110100011100, 
24'b001001111001001011101011, 
24'b110101011111110100010010, 
24'b001011000111001011101110, 
24'b110100011001110100010101, 
24'b001100000001001011100101, 
24'b110011101011110100100010, 
24'b001100100000001011010010, 
24'b110011011100110100111101, 
24'b001100100000001010110001, 
24'b110011101110110101100110, 
24'b001011111100001001111111, 
24'b110100100011110110100000, 
24'b001010111000001000111100, 
24'b110101110110110111101100, 
24'b001001010101000111100110, 
24'b110111100101111001001100, 
24'b000111011100000101111011, 
24'b111001100110111010111111, 
24'b000101010100000100000001, 
24'b111011110001111101000011, 
24'b000011001011000001110110, 
24'b111101111000111111010010, 
24'b000001001010111111100100, 
24'b111111101111000001100111, 
24'b111111011101111101001110, 
24'b000001001110000011111010, 
24'b111110010001111011000001, 
24'b000010000111000110000010, 
24'b111101101101111001000001, 
24'b000010010101000111110111, 
24'b111101110111110111011010, 
24'b000001110010001001001110, 
24'b111110110001110110010010, 
24'b000000100000001010000100, 
24'b000000011010110101101111, 
24'b111110100010001010010101, 
24'b000010101100110101110011, 
24'b111011111111001001111011, 
24'b000101011110110110100000, 
24'b111001000010001000111100, 
24'b001000100010110111110010, 
24'b110101111010000111011000, 
24'b001011101010111001100010, 
24'b110010110101000101011110, 
24'b001110100101111011101000, 
24'b110000000110000011010010, 
24'b010001000101111101111000, 
24'b101101111010000001000000, 
24'b010010111001000000000110, 
24'b101100100000111110111000, 
24'b010011111000000010000111, 
24'b101100000000111101000000, 
24'b010011111000000011110000, 
24'b101100100011111011101000, 
24'b010010110100000100111000, 
24'b101110000101111010110001, 
24'b010000110001000101011010, 
24'b110000100110111010100100, 
24'b001101110100000101010110, 
24'b110011111101111010111100, 
24'b001010000111000100101001, 
24'b110111111101111011111010, 
24'b000101111010000011011110, 
24'b111100010100111101010001, 
24'b000001011101000001111100, 
24'b000000110001111110111011, 
24'b111101000101000000001110, 
24'b000101000001000000101010, 
24'b111001000010111110100000, 
24'b001000110010000010010010, 
24'b110101100110111101000010, 
24'b001011110101000011100101, 
24'b110010111111111011111100, 
24'b001101111110000100011010, 
24'b110001010100111011011010, 
24'b001111001001000100101000, 
24'b1_10000101010111011100010,
24'b000101100110000001110111, 
24'b111011000001111110001101, 
24'b000100010111000001101110, 
24'b111100010010111110010110, 
24'b000011000100000001100111, 
24'b111101101000111110011101, 
24'b000001101101000001100000, 
24'b111110111110111110100010, 
24'b000000010110000001011011, 
24'b000000010101111110100111, 
24'b111111000001000001011001, 
24'b000001101000111110100111, 
24'b111101101111000001011001, 
24'b000010111001111110100111, 
24'b111100100000000001011011, 
24'b000100000011111110100011, 
24'b111011011010000001100000, 
24'b000101000111111110011101, 
24'b111010011010000001100110, 
24'b000110000010111110010101, 
24'b111001100101000001110000, 
24'b000110110010111110001100, 
24'b111000111010000001111011, 
24'b000111010110111110000000, 
24'b111000011011000010000101, 
24'b000111110001111101110101, 
24'b111000000111000010010010, 
24'b000111111110111101100111, 
24'b110111111111000010011110, 
24'b001000000000111101011100, 
24'b111000000011000010101010, 
24'b000111110110111101010001, 
24'b111000010001000010110100, 
24'b000111100100111101001000, 
24'b111000101011000010111100, 
24'b000111000100111101000001, 
24'b111001001111000011000010, 
24'b000110011101111100111100, 
24'b111001111010000011000101, 
24'b000101101101111100111011, 
24'b111010101100000011000100, 
24'b000100111001111100111101, 
24'b111011100011000011000010, 
24'b000011111111111101000010, 
24'b111100011111000010111010, 
24'b000011000100111101001011, 
24'b111101011010000010101111, 
24'b000010000111111101010111, 
24'b111110010110000010100001, 
24'b000001001101111101100111, 
24'b111111001111000010001111, 
24'b000000010101111101111010, 
24'b000000000100000001111011, 
24'b111111100011111110010000, 
24'b000000110011000001100100, 
24'b111110110111111110101000, 
24'b000001011011000001001011, 
24'b111110010011111111000010, 
24'b000001111011000000110001, 
24'b111101111000111111011101, 
24'b000010010010000000010110, 
24'b111101100110111111110111, 
24'b000010011110111111111011, 
24'b111101011111000000010001, 
24'b000010100000111111100011, 
24'b111101100010000000101001, 
24'b000010011000111111001100, 
24'b111101110000000000111111, 
24'b000010000110111110110110, 
24'b111110000111000001010011, 
24'b000001101010111110100101, 
24'b111110100111000001100010, 
24'b000001000110111110011000, 
24'b111111001111000001101110, 
24'b000000011010111110001110, 
24'b111111111110000001110100, 
24'b111111101000111110001010, 
24'b000000110001000001110110, 
24'b111110110010111110001010, 
24'b000001101010000001110100, 
24'b111101111010111110001111, 
24'b000010100010000001101100, 
24'b111101000000111110011010, 
24'b000011011011000001100000, 
24'b111100001010111110101000, 
24'b000100010001000001001111, 
24'b111011010101111110111011, 
24'b000101000011000000111010, 
24'b111010100110111111010001, 
24'b000101101111000000100010, 
24'b111001111101111111101010, 
24'b000110010010000000001000, 
24'b111001011111000000000110, 
24'b000110101101111111101100, 
24'b111001001001000000100010, 
24'b000110111100111111010000, 
24'b111001000000000000111110, 
24'b000110111111111110110100, 
24'b111001000011000001011001, 
24'b000110110111111110011010, 
24'b111001010011000001110010, 
24'b000110100000111110000011, 
24'b111001101111000010000111, 
24'b000101111110111101110000, 
24'b111010011001000010011000, 
24'b000101001110111101100011, 
24'b111011001111000010100010, 
24'b000100010001111101011010, 
24'b111100010010000010100111, 
24'b000011001010111101011001, 
24'b111101011110000010100101, 
24'b000001111001111101100000, 
24'b111110110011000010011011, 
24'b000000100000111101101110, 
24'b000000010000000010001000, 
24'b111111000000111110000101, 
24'b000001110010000001101100, 
24'b111101011011111110100101, 
24'b000011011000000001001001, 
24'b111011110101111111001100, 
24'b000100111111000000011101, 
24'b111010001110111111111100, 
24'b000110100100111111101001, 
24'b111000101010000000110011, 
24'b001000000111111110101110, 
24'b110111001011000001110010, 
24'b001001100010111101101101, 
24'b110101110010000010110110, 
24'b001010110111111100100110, 
24'b110100100010000011111111, 
24'b001100000010111011011011, 
24'b110011011101000101001011, 
24'b001101000001111010001101, 
24'b110010100100000110011001, 
24'b001101110011111000111111, 
24'b110001111010000111101000, 
24'b001110010111110111110001, 
24'b110001011100001000110101, 
24'b001110101100110110100101, 
24'b110001001111001010000000, 
24'b001110110010110101011101, 
24'b110001010001001011000110, 
24'b001110101000110100011010, 
24'b110001100011001100000101, 
24'b001110001111110011011110, 
24'b110010000011001100111101, 
24'b001101101000110010101010, 
24'b110010110000001101101100, 
24'b001100110101110001111111, 
24'b110011101010001110010001, 
24'b001011110100110001100000, 
24'b110100101111001110101011, 
24'b001010101011110001001101, 
24'b110101111100001110111000, 
24'b001001011001110001000101, 
24'b110111010010001110111001, 
24'b001000000001110001001100, 
24'b111000101011001110101100, 
24'b000110100111110001011110, 
24'b111010001000001110010010, 
24'b000101001011110010000000, 
24'b111011100011001101101100, 
24'b000011110000110010101101, 
24'b111100111011001100110111, 
24'b000010011011110011100111, 
24'b111110001110001011110111, 
24'b000001001011110100101100, 
24'b111111011010001010101100, 
24'b000000000011110101111110, 
24'b000000011100001001010110, 
24'b111111000110110111010111, 
24'b000001010100000111111000, 
24'b111110010101111000111001, 
24'b000001111101000110010010, 
24'b111101110010111010100010, 
24'b000010011010000100100111, 
24'b111101011110111100010000, 
24'b000010100110000010111000, 
24'b111101011001111101111111, 
24'b000010100011000001001000, 
24'b111101100100111111110001, 
24'b000010010000111111010110, 
24'b111101111111000001100010, 
24'b000001101111111101100110, 
24'b111110100111000011010001, 
24'b000000111110111011111001, 
24'b111111011110000100111011, 
24'b000000000010111010010001, 
24'b000000100001000110100000, 
24'b111110111000111000110000, 
24'b000001110000000111111110, 
24'b111101100101110111010110, 
24'b000011000111001001010011, 
24'b111100001010110110000110, 
24'b000100100101001010011111, 
24'b111010101010110100111111, 
24'b000110000111001011100001, 
24'b111001000110110100000010, 
24'b000111101100001100010111, 
24'b110111100010110011010010, 
24'b001001001111001101000010, 
24'b110110000001110010101101, 
24'b001010101111001101100001, 
24'b110100100100110010010100, 
24'b001100000111001101110011, 
24'b110011001111110010000111, 
24'b001101011001001101111100, 
24'b110010000011110010000101, 
24'b001110011111001101111000, 
24'b110001000011110010001110, 
24'b001111011000001101101001, 
24'b110000010000110010100001, 
24'b010000000011001101010001, 
24'b101111101110110010111110, 
24'b010000011110001100110000, 
24'b101111011100110011100011, 
24'b010000100110001100000111, 
24'b101111011011110100001111, 
24'b010000011111001011011000, 
24'b101111101101110101000010, 
24'b010000000100001010100011, 
24'b110000010000110101111001, 
24'b001111011000001001101010, 
24'b110001000101110110110100, 
24'b001110011010001000101101, 
24'b110010001010110111110001, 
24'b001101001101000111110000, 
24'b110011011111111000110000, 
24'b001011110001000110110000, 
24'b110101000010111001101110, 
24'b001010000111000101110010, 
24'b110110110001111010101101, 
24'b001000010011000100110101, 
24'b111000101010111011101001, 
24'b000110010110000011111011, 
24'b111010101011111100100010, 
24'b000100010010000011000011, 
24'b111100110000111101011000, 
24'b000010001011000010001111, 
24'b111110111010111110001010, 
24'b000000000011000001011111, 
24'b000001000001111110110111, 
24'b111101111100000000110011, 
24'b000011000110111111100001, 
24'b111011111000000000001100, 
24'b000101000110000000000110, 
24'b111001111100111111101011, 
24'b000110111110000000100100, 
24'b111000001001111111001110, 
24'b001000101011000000111110, 
24'b110110100010111110110101, 
24'b001010001110000001010101, 
24'b110101000110111110100011, 
24'b001011100001000001100110, 
24'b110011111010111110010100, 
24'b001100100111000001110011, 
24'b110010111101111110001001, 
24'b001101011011000001111100, 
24'b110010010001111110000001, 
24'b001101111111000010000001, 
24'b110001110110111101111111, 
24'b001110010010000010000011, 
24'b110001101010111101111110, 
24'b001110010101000010000001, 
24'b110001110001111110000001, 
24'b001110000111000001111101, 
24'b110010000110111110000111, 
24'b001101101001000001110101, 
24'b110010101011111110001111, 
24'b001100111110000001101100, 
24'b110011011100111110011010, 
24'b001100000111000001011111, 
24'b110100011010111110100111, 
24'b001011000100000001010011, 
24'b110101100000111110110101, 
24'b001001111001000001000010, 
24'b110110101110111111000111, 
24'b001000101000000000110000, 
24'b111000000001111111011010, 
24'b000111010100000000011010, 
24'b111001011000111111110001, 
24'b000101111101000000000100, 
24'b111010110000000000001001, 
24'b000100100101111111101010, 
24'b111100000100000000100100, 
24'b000011010011111111001110, 
24'b111101010110000001000011, 
24'b000010000100111110101101, 
24'b111110100001000001100100, 
24'b000000111101111110001100, 
24'b111111100101000010001000, 
24'b111111111110111101100100, 
24'b000000011110000010110000, 
24'b111111001001111100111011, 
24'b000001001101000011011010, 
24'b111110100001111100001110, 
24'b000001101111000100001010, 
24'b111110000100111011011110, 
24'b000010000101000100111100, 
24'b111101110101111010101011, 
24'b000010001101000101110000, 
24'b111101110100111001110100, 
24'b000010001001000110101001, 
24'b111101111111111000111010, 
24'b000001110110000111100100, 
24'b111110011000110111111111, 
24'b000001011001001000100000, 
24'b111110111100110111000000, 
24'b000000101110001001011111, 
24'b111111101100110110000001, 
24'b111111111000001010100000, 
24'b000000100111110101000000, 
24'b111110111000001011100000, 
24'b000001101001110011111111, 
24'b111101110010001100100000, 
24'b000010110100110011000000, 
24'b111100100101001101011111, 
24'b000100000011110010000010, 
24'b111011010101001110011100, 
24'b000101010101110001000110, 
24'b111010000010001111010111, 
24'b000110101001110000001101, 
24'b111000101101010000001110, 
24'b000111111101101111011000, 
24'b110111011010010000111111, 
24'b001001001110101110101001, 
24'b110110001010010001101101, 
24'b001010011100101101111111, 
24'b110100111111010010010100, 
24'b001011100100101101011011, 
24'b110011111010010010110100, 
24'b001100100110101100111111, 
24'b110010111100010011001100, 
24'b001101011111101100101011, 
24'b110010001000010011011011, 
24'b001110001111101100100000, 
24'b110001011100010011100011, 
24'b001110110110101100011100, 
24'b110000111011010011100001, 
24'b001111010010101100100010, 
24'b110000100100010011010111, 
24'b001111100100101100110010, 
24'b110000010111010011000011, 
24'b001111101011101101001010, 
24'b110000010110010010101000, 
24'b001111101001101101101010, 
24'b110000011101010010000010, 
24'b001111011011101110010011, 
24'b110000101111010001010101, 
24'b001111000110101111000101, 
24'b110001001001010000011111, 
24'b001110100111101111111110, 
24'b110001101001001111100011, 
24'b001110000011110000111110, 
24'b110010010001001110100000, 
24'b001101011001110010000100, 
24'b110010111101001101010110, 
24'b001100101010110011010000, 
24'b110011101111001100001001, 
24'b001011111001110100011111, 
24'b110100100000001010111000, 
24'b001011000110110101110010, 
24'b110101010100001001100011, 
24'b001010010011110111001000, 
24'b110110000111001000001100, 
24'b001001100001111000011111, 
24'b110110111001000110110101, 
24'b001000110001111001110111, 
24'b110111100110000101011100, 
24'b001000000100111011001110, 
24'b111000010000000100000110, 
24'b000111011100111100100100, 
24'b111000110111000010110001, 
24'b000110111010111101111001, 
24'b111001010110000001011101, 
24'b000110011100111111001010, 
24'b111001110000000000001111, 
24'b000110000101000000010111, 
24'b111010000100111111000011, 
24'b000101110101000001100001, 
24'b111010010010111101111100, 
24'b000101101011000010100110, 
24'b111010011001111100111010, 
24'b000101100110000011100101, 
24'b111010011010111011111101, 
24'b000101101000000100011111, 
24'b111010010111111011000101, 
24'b000101101101000101010100, 
24'b111010001111111010010100, 
24'b000101110111000110000011, 
24'b111010000010111001101000, 
24'b000110000101000110101100, 
24'b111001110011111001000011, 
24'b000110010100000111001110, 
24'b111001100011111000100011, 
24'b000110100101000111101011, 
24'b111001010010111000001001, 
24'b000110110111001000000010, 
24'b111001000010110111110100, 
24'b000111000110001000010011, 
24'b111000110100110111100110, 
24'b000111010011001000011110, 
24'b111000101000110111011101, 
24'b000111011100001000100110, 
24'b111000100001110111011000, 
24'b000111100001001000100111, 
24'b111000011111110111011011, 
24'b000111011111001000100011, 
24'b111000100100110111100001, 
24'b000111010111001000011010, 
24'b111000101110110111101100, 
24'b000111001000001000001101, 
24'b111001000010110111111011, 
24'b000110110011000111111100, 
24'b111001011011111000001111, 
24'b000110010100000111100110, 
24'b111001111101111000100111, 
24'b000101101110000111001011, 
24'b111010101000111001000011, 
24'b000101000000000110101101, 
24'b111011011011111001100010, 
24'b000100001010000110001100, 
24'b111100010100111010000111, 
24'b000011001100000101100111, 
24'b111101010110111010101101, 
24'b000010001000000100111110, 
24'b111110011100111011011000, 
24'b000000111110000100010011, 
24'b111111101001111100000100, 
24'b111111110001000011100011, 
24'b000000110111111100110101, 
24'b111110011111000010110011, 
24'b000010001010111101100111, 
24'b111101001101000001111111, 
24'b000011011110111110011100, 
24'b111011111000000001001001, 
24'b000100110001111111010010, 
24'b111010100101000000010010, 
24'b000110000011000000001010, 
24'b111001010101111111011010, 
24'b000111010011000001000010, 
24'b111000001001111110100001, 
24'b001000011100000001111011, 
24'b110111000001111101101001, 
24'b001001100000000010110011, 
24'b110110000010111100110010, 
24'b001010011011000011101001, 
24'b110101001001111011111100, 
24'b001011001111000100011110, 
24'b110100011011111011001001, 
24'b001011111000000101010000, 
24'b110011111000111010010111, 
24'b001100010101000101111111, 
24'b110011100001111001101011, 
24'b001100101000000110101010, 
24'b110011010100111001000011, 
24'b001100101101000111010000, 
24'b110011010110111000011111, 
24'b001100100101000111110001, 
24'b110011100100111000000001, 
24'b001100001111001000001100, 
24'b110100000000110111101010, 
24'b001011101100001000011111, 
24'b110100101010110111011001, 
24'b001010111101001000101100, 
24'b110101011111110111010000, 
24'b001010000000001000110010, 
24'b110110100010110111001101, 
24'b001000110111001000110001, 
24'b110111110010110111010011, 
24'b000111100100001000101000, 
24'b111001001010110111011111, 
24'b000110000101001000011001, 
24'b111010101101110111110010, 
24'b000100011111001000000001, 
24'b111100010111111000001100, 
24'b000010110010000111100110, 
24'b111110000111111000101011, 
24'b000000111110000111000011, 
24'b111111111101111001010000, 
24'b111111000111000110011100, 
24'b000001110101111001111010, 
24'b111101001101000101110001, 
24'b000011110000111010100110, 
24'b111011010100000101000011, 
24'b000101101001111011010100, 
24'b111001011100000100010100, 
24'b000111100000111100000100, 
24'b110111101000000011100101, 
24'b001001010000111100110010, 
24'b110101111001000010110111, 
24'b001010111101111101100000, 
24'b110100010010000010001100, 
24'b001100011101111110001001, 
24'b110010110100000001100101, 
24'b001101111000111110101110, 
24'b110001100001000001000010, 
24'b001111000100111111001100, 
24'b110000011001000000100111, 
24'b010000000110111111100100, 
24'b101111011111000000010100, 
24'b010000111001111111110010, 
24'b101110110101000000001010, 
24'b010001011100111111110111, 
24'b101110011010000000001010, 
24'b010001101111111111110001, 
24'b101110001110000000010100, 
24'b010001110010111111100010, 
24'b101110010011000000101011, 
24'b010001100100111111000110, 
24'b101110101001000001001011, 
24'b010001000111111110100000, 
24'b101111001111000001110111, 
24'b010000011000111101101111, 
24'b110000000110000010101111, 
24'b001111011001111100110010, 
24'b110001001101000011110000, 
24'b001110001010111011101011, 
24'b110010100010000100111011, 
24'b001100101101111010011100, 
24'b110100000111000110001111, 
24'b001011000011111001000101, 
24'b110101111000000111101010, 
24'b001001001100110111100111, 
24'b110111110100001001001001, 
24'b000111001011110110000111, 
24'b111001111010001010101101, 
24'b000101000000110100100010, 
24'b111100000111001100010001, 
24'b000010101111110010111100, 
24'b111110011100001101110111, 
24'b000000010111110001011000, 
24'b000000110110001111011001, 
24'b111101111101101111111001, 
24'b000011010010010000110111, 
24'b111011100000101110011101, 
24'b000101101110010010001101, 
24'b111001000101101101001011, 
24'b001000001010010011011011, 
24'b110110101011101100000011, 
24'b001010100001010100011101, 
24'b110100010101101011000111, 
24'b001100110100010101010011, 
24'b110010000100101010011000, 
24'b001111000000010101111010, 
24'b101111111100101001111001, 
24'b010001000110010110010010, 
24'b101101111100101001101001, 
24'b010011000001010110011001, 
24'b101100000110101001101011, 
24'b010100110001010110001110, 
24'b101010011010101001111110, 
24'b010110010110010101110001, 
24'b101000111100101010100101, 
24'b010111101111010101000011, 
24'b100111101001101011011100, 
24'b011000111010010100000010, 
24'b100110100101101100100101, 
24'b011001110111010010110001, 
24'b100101101110101101111111, 
24'b011010101001010001001111, 
24'b100101000101101111101000, 
24'b011011001100001111011111, 
24'b100100100111110001011110, 
24'b011011100011001101100001, 
24'b100100010111110011100010, 
24'b011011101101001011011010, 
24'b100100010011110101101101, 
24'b011011101011001001001001, 
24'b100100011010111000000001, 
24'b011011011110000110110011, 
24'b100100101100111010011010, 
24'b011011001000000100011000, 
24'b100101000110111100110110, 
24'b011010101000000001111101, 
24'b100101101010111111010000, 
24'b011010000010111111100011, 
24'b100110010101000001101000, 
24'b011001010011111101001110, 
24'b100111000101000011111011, 
24'b011000100001111010111111, 
24'b100111111001000110000100, 
24'b010111101011111000111010, 
24'b101000110001001000000100, 
24'b010110110010110111000001, 
24'b101001101011001001110110, 
24'b010101110111110101010110, 
24'b101010100110001011011010, 
24'b010100111110110011111010, 
24'b101011011111001100101101, 
24'b010100000010110010101111, 
24'b101100011010001101101111, 
24'b010011001010110001110110, 
24'b101101010010001110011111, 
24'b010010010010110001010000, 
24'b101110001000001110111100, 
24'b010001011110110000111100, 
24'b101110111011001111000101, 
24'b010000101101110000111101, 
24'b101111101011001110111101, 
24'b001111111110110001001110, 
24'b110000011000001110100010, 
24'b001111010001110001110010, 
24'b110001000010001101110110, 
24'b001110101001110010100110, 
24'b110001101001001100111001, 
24'b001110000010110011101001, 
24'b110010001111001011110001, 
24'b001101011111110100111000, 
24'b110010110010001010011011, 
24'b001100111011110110010100, 
24'b110011010110001000111100, 
24'b001100011010110111110110, 
24'b110011110111000111010110, 
24'b001011110111111001100001, 
24'b110100011010000101101011, 
24'b001011010100111011001100, 
24'b110100111110000011111101, 
24'b001010110000111100111010, 
24'b110101100011000010010000, 
24'b001010001000111110100101, 
24'b110110001100000000100110, 
24'b001001011110000000001101, 
24'b110110111000111111000011, 
24'b001000110001000001101110, 
24'b110111100111111101100100, 
24'b000111111111000011000111, 
24'b111000011100111100010001, 
24'b000111001000000100010101, 
24'b111001010110111011001001, 
24'b000110001011000101010111, 
24'b111010010100111010001101, 
24'b000101001010000110001011, 
24'b111011011001111001100000, 
24'b000100000100000110110010, 
24'b111100100000111001000001, 
24'b000010111000000111001000, 
24'b111101101111111000110010, 
24'b000001101000000111010000, 
24'b111111000010111000110010, 
24'b000000010100000111001000, 
24'b000000010110111001000001, 
24'b111110111101000110110010, 
24'b000001101111111001011110, 
24'b111101100100000110001111, 
24'b000011001010111010001001, 
24'b111100001001000101011101, 
24'b000100100101111011000000, 
24'b111010101110000100100001, 
24'b000101111111111100000001, 
24'b111001010100000011011100, 
24'b000111010111111101001010, 
24'b110111111101000010001110, 
24'b001000101101111110011011, 
24'b110110101010000000111010, 
24'b001001111101111111110001, 
24'b110101011100111111100010, 
24'b001011001001000001001010, 
24'b110100010101111110001010, 
24'b001100001101000010100010, 
24'b110011010101111100110010, 
24'b001101001000000011111001, 
24'b110010011110111011011100, 
24'b001101111010000101001101, 
24'b110001110001111010001101, 
24'b001110100010000110011010, 
24'b110001001110111001000011, 
24'b001110111111000111011111, 
24'b110000110111111000000001, 
24'b001111001111001000011010, 
24'b110000101100110111001011, 
24'b001111010101001001001101, 
24'b110000101100110110011111, 
24'b001111001110001001110010, 
24'b110000111001110101111110, 
24'b001110111101001010001100, 
24'b110001010000110101101011, 
24'b001110100000001010011000, 
24'b110001110011110101100101, 
24'b001101111000001010011001, 
24'b110010011111110101101100, 
24'b001101000111001010001011, 
24'b110011010110110101111111, 
24'b001100001110001001110010, 
24'b110100010010110110100000, 
24'b001011001011001001001100, 
24'b110101010111110111001011, 
24'b001010000110001000011100, 
24'b110110011111110111111111, 
24'b001000111011000111100011, 
24'b110111101011111000111101, 
24'b000111101110000110100001, 
24'b111000111000111010000010, 
24'b000110100000000101011010, 
24'b111010000110111011001101, 
24'b000101010101000100001101, 
24'b111011010000111100011010, 
24'b000100001100000010111110, 
24'b111100010111111101101001, 
24'b000011000111000001101111, 
24'b111101011000111110111001, 
24'b000010001010000000100000, 
24'b111110010011000000000111, 
24'b000001010100111111010101, 
24'b111111000100000001001111, 
24'b000000100101111110001101, 
24'b111111101101000010010011, 
24'b000000000010111101001110, 
24'b000000001100000011010000, 
24'b111111101001111100010101, 
24'b000000011111000100000011, 
24'b111111011101111011100111, 
24'b000000100110000100101101, 
24'b111111011011111011000010, 
24'b000000100010000101001100, 
24'b111111100100111010101001, 
24'b000000010011000101011111, 
24'b111111111001111010011100, 
24'b111111111001000101100110, 
24'b000000010111111010011100, 
24'b111111010101000101100000, 
24'b000001000000111010100111, 
24'b111110101000000101001110, 
24'b000001110010111011000000, 
24'b111101110011000100110000, 
24'b000010101001111011100100, 
24'b111100111000000100000110, 
24'b000011101000111100010011, 
24'b111011111000000011010001, 
24'b000100101001111101001101, 
24'b111010110100000010010010, 
24'b000101101101111110010001, 
24'b111001110000000001001010, 
24'b000110110001111111011110, 
24'b111000101101111111111010, 
24'b000111110100000000110000, 
24'b110111101100111110100101, 
24'b001000110011000010001000, 
24'b110110101111111101001001, 
24'b001001101101000011100101, 
24'b110101111000111011101101, 
24'b001010100001000101000010, 
24'b110101001000111010001110, 
24'b001011001100000110100010, 
24'b110100100010111000101111, 
24'b001011101110000111111111, 
24'b110100000101110111010011, 
24'b001100000101001001011011, 
24'b110011110011110101111001, 
24'b001100010001001010110001, 
24'b110011101110110100100101, 
24'b001100010001001100000011, 
24'b110011110011110011010111, 
24'b001100000101001101001101, 
24'b110100000101110010010001, 
24'b001011101110001110001111, 
24'b110100100010110001010100, 
24'b001011001011001111000111, 
24'b110101001011110000100001, 
24'b001010011101001111110110, 
24'b110101111110101111111000, 
24'b001001100101010000011000, 
24'b110110111011101111011100, 
24'b001000100100010000101110, 
24'b110111111111101111001011, 
24'b000111011100010000111001, 
24'b111001001010101111000111, 
24'b000110001111010000110111, 
24'b111010011010101111001111, 
24'b000100111101010000101000, 
24'b111011101110101111100100, 
24'b000011101000010000001110, 
24'b111101000011110000000110, 
24'b000010010011001111100110, 
24'b111110010111110000110011, 
24'b000001000000001110110011, 
24'b111111101000110001101100, 
24'b111111110000001101110011, 
24'b000000110110110010110001, 
24'b111110100110001100101010, 
24'b000001111110110011111111, 
24'b111101100010001011010111, 
24'b000010111111110101011000, 
24'b111100100101001001111001, 
24'b000011110110110110110111, 
24'b111011110010001000010110, 
24'b000100100101111000011111, 
24'b111011001001000110101100, 
24'b000101001000111010001101, 
24'b111010101011000100111011, 
24'b000101100001111100000000, 
24'b111010010111000011000101, 
24'b000101101101111101110110, 
24'b111010010001000001001110, 
24'b000101101111111111101111, 
24'b111010010110111111010101, 
24'b000101100100000001100111, 
24'b111010100101111101011100, 
24'b000101001111000011100001, 
24'b111011000000111011100100, 
24'b000100110000000101010111, 
24'b111011100100111001101111, 
24'b000100001000000111001010, 
24'b111100010000110111111110, 
24'b000011010110001000111000, 
24'b111101000100110110010100, 
24'b000010100000001010100001, 
24'b111101111110110100101110, 
24'b000001100100001100000001, 
24'b111110111100110011010010, 
24'b000000100100001101011001, 
24'b111111111101110001111111, 
24'b111111100010001110100110, 
24'b000000111111110000110111, 
24'b111110100001001111101001, 
24'b000010000001101111111010, 
24'b111101011111010000011111, 
24'b000011000001101111001011, 
24'b111100100001010001001000, 
24'b000011111101101110101000, 
24'b111011100110010001100100, 
24'b000100110100101110010011, 
24'b111010110010010001110001, 
24'b000101100111101110001101, 
24'b111010000100010001110001, 
24'b000110010001101110010110, 
24'b111001011101010001100001, 
24'b000110110101101110101101, 
24'b111000111101010001000001, 
24'b000111010000101111010011, 
24'b111000100110010000010011, 
24'b000111100100110000001001, 
24'b111000010110001111010111, 
24'b000111101110110001001101, 
24'b111000001111001110001011, 
24'b000111110001110010011111, 
24'b111000001111001100110100, 
24'b000111101100110011111100, 
24'b111000011001001011010000, 
24'b000111100001110101100111, 
24'b111000101000001001100000, 
24'b000111001110110111011011, 
24'b111000111101000111100110, 
24'b000110111000111001011010, 
24'b111001010101000101100100, 
24'b000110011100111011011111, 
24'b111001110010000011011011, 
24'b000101111111111101101100, 
24'b111010010001000001001100, 
24'b000101011110111111111011, 
24'b111010110010111110111011, 
24'b000100111111000010001111, 
24'b111011010001111100101000, 
24'b000100011111000100100010, 
24'b111011110000111010010101, 
24'b000100000010000110110100, 
24'b111100001100111000000101, 
24'b000011100111001001000010, 
24'b111100100101110101111001, 
24'b000011010001001011001011, 
24'b111100111010110011110011, 
24'b000010111110001101001100, 
24'b111101001001110001110110, 
24'b000010110000001111000100, 
24'b111101010101110000000011, 
24'b000010101000010000110010, 
24'b111101011010101110011100, 
24'b000010100110010010010011, 
24'b111101011010101101000001, 
24'b000010101000010011100111, 
24'b111101010110101011110101, 
24'b000010101111010100101101, 
24'b111101001011101010110110, 
24'b000010111011010101100011, 
24'b111100111101101010001001, 
24'b000011001100010110001000, 
24'b111100101100101001101011, 
24'b000011011111010110011101, 
24'b111100010111101001011110, 
24'b000011110100010110100010, 
24'b111100000001101001100010, 
24'b000100001010010110010111, 
24'b111011101010101001110100, 
24'b000100100001010101111101, 
24'b111011010101101010010111, 
24'b000100110110010101010011, 
24'b111011000000101011000111, 
24'b000101001001010100011100, 
24'b111010110000101100000100, 
24'b000101011001010011011010, 
24'b111010100010101101001100, 
24'b000101100011010010001100, 
24'b111010011001101110011111, 
24'b000101101001010000110100, 
24'b111010010111101111111010, 
24'b000101101001001111010111, 
24'b111010011010110001011011, 
24'b000101100010001101110011, 
24'b111010100101110010111111, 
24'b000101010011001100001110, 
24'b111010110110110100100111, 
24'b000100111111001010100110, 
24'b111011001111110110001101, 
24'b000100100010001001000001, 
24'b111011110000110111110001, 
24'b000011111110000111011111, 
24'b111100010110111001010001, 
24'b000011010100000110000010, 
24'b111101000100111010101011, 
24'b000010100101000100101011, 
24'b111101110101111011111101, 
24'b000001110000000011011110, 
24'b111110101100111101000110, 
24'b000000111000000010011010, 
24'b111111100110111110000100, 
24'b111111111100000001100010, 
24'b000000100001111110110101, 
24'b111111000001000000110110, 
24'b000001011110111111011100, 
24'b111110000100000000010110, 
24'b000010011011111111110100, 
24'b111101001000000000000101, 
24'b000011010100111111111111, 
24'b111100010001000000000000, 
24'b000100001011111111111101, 
24'b111011011011000000001000, 
24'b000100111101111111101110, 
24'b111010101101000000011101, 
24'b000101101001111111010100, 
24'b111010000100000000111101, 
24'b000110001110111110101110, 
24'b111001100010000001101001, 
24'b000110101100111101111110, 
24'b111001001000000010011110, 
24'b000111000010111101000101, 
24'b111000111000000011011011, 
24'b000111001110111100000100, 
24'b111000101110000100011111, 
24'b000111010010111010111110, 
24'b111000110000000101100111, 
24'b000111001101111001110100, 
24'b111000111001000110110000, 
24'b000111000000111000101001, 
24'b111001001010000111111101, 
24'b000110101010110111011101, 
24'b111001100100001001001000, 
24'b000110001110110110010100, 
24'b111010000011001010010000, 
24'b000101101010110101001101, 
24'b111010101001001011010011, 
24'b000101000010110100001100, 
24'b111011010011001100010010, 
24'b000100010111110011010001, 
24'b111100000000001101001001, 
24'b000011101001110010011111, 
24'b111100101111001101110111, 
24'b000010111001110001110101, 
24'b111101011110001110011100, 
24'b000010001100110001010101, 
24'b111110001011001110110111, 
24'b000001011111110001000000, 
24'b111110110101001111000111, 
24'b000000111000110000110101, 
24'b111111011011001111001100, 
24'b000000010100110000110110, 
24'b111111111011001111000101, 
24'b111111111000110001000001, 
24'b000000010100001110110100, 
24'b111111100010110001011000, 
24'b000000100110001110011001, 
24'b111111010101110001110111, 
24'b000000101111001101110100, 
24'b111111010000110010100001, 
24'b000000101111001101000110, 
24'b111111010101110011010011, 
24'b000000100100001100010001, 
24'b111111100011110100001100, 
24'b000000010011001011010101, 
24'b111111111010110101001011, 
24'b111111110111001010010101, 
24'b000000011010110110001111, 
24'b111111010011001001001111, 
24'b000001000001110111010101, 
24'b111110101000001000001000, 
24'b000001110000111000011100, 
24'b111101110111000110111111, 
24'b000010100100111001100101, 
24'b111101000000000101110111, 
24'b000011011101111010101101, 
24'b111100000110000100110000, 
24'b000100011000111011110010, 
24'b111011001010000011101100, 
24'b000101010101111100110101, 
24'b111010001101000010101100, 
24'b000110010001111101110001, 
24'b111001010011000001110001, 
24'b000111001010111110101011, 
24'b111000011011000000111011, 
24'b001000000000111111011110, 
24'b110111100111000000001011, 
24'b001000110000000000001011, 
24'b110110111011111111100001, 
24'b001001011000000000110000, 
24'b110110010110111110111111, 
24'b001001111001000001010001, 
24'b110101111011111110100010, 
24'b001010001110000001101001, 
24'b110101101010111110001100, 
24'b001010011010000001111100, 
24'b110101100101111101111101, 
24'b001010011010000010001001, 
24'b110101101011111101110010, 
24'b001010001111000010010001, 
24'b110101111100111101101110, 
24'b001001111000000010010011, 
24'b110110011000111101101100, 
24'b001001010100000010010011, 
24'b110111000001111101110000, 
24'b001000100111000010001110, 
24'b110111110100111101110101, 
24'b000111110000000010001000, 
24'b111000110000111101111100, 
24'b000110101110000010000000, 
24'b111001110101111110000101};