logic [23:0] sig_pr [0:2047] = {
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111110000000000101,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111110000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000101,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b111111111111000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000110,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000000000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000001000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000000111,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000010000000001000,
24'b111111111111000000000000,
24'b000000000011000000000111,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000011000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001000,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000100000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000101000000001001,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001001,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000110000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000000111000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001010000000001011,
24'b000000000000000000000000,
24'b000000001010000000001011,
24'b000000000000000000000000,
24'b000000001010000000001011,
24'b000000000000000000000000,
24'b000000001010000000001100,
24'b000000000000000000000000,
24'b000000001010000000001100,
24'b000000000000000000000000,
24'b000000001010000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001011000000001100,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001101,
24'b000000000000000000000000,
24'b000000001100000000001100,
24'b000000000000000000000000,
24'b000000001100000000001101,
24'b000000000000000000000000,
24'b000000001100000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001101000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001110000000001101,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000001111000000001110,
24'b000000000000000000000000,
24'b000000010000000000001110,
24'b000000000000000000000000,
24'b000000010000000000001110,
24'b000000000000000000000000,
24'b000000010000000000001110,
24'b000000000000000000000000,
24'b000000010001000000001110,
24'b000000000000000000000000,
24'b000000010001000000001110,
24'b000000000000000000000000,
24'b000000010001000000001111,
24'b000000000000000000000000,
24'b000000010001000000001111,
24'b000000000000000000000000,
24'b000000010010000000001111,
24'b000000000000000000000000,
24'b000000010010000000001111,
24'b000000000000000000000000,
24'b000000010010000000001111,
24'b000000000000000000000000,
24'b000000010011000000001111,
24'b000000000000000000000000,
24'b000000010011000000001111,
24'b000000000000000000000000,
24'b000000010011000000001111,
24'b000000000000000000000000,
24'b000000010100000000010000,
24'b000000000000000000000000,
24'b000000010100000000010000,
24'b000000000000000000000000,
24'b000000010100000000010000,
24'b000000000000000000000000,
24'b000000010101000000010000,
24'b000000000000000000000000,
24'b000000010101000000010000,
24'b000000000000000000000000,
24'b000000010110000000010000,
24'b000000000000000000000000,
24'b000000010110000000010000,
24'b000000000000000000000000,
24'b000000010110000000010000,
24'b000000000000000000000000,
24'b000000010111000000010001,
24'b000000000000000000000000,
24'b000000010111000000010001,
24'b000000000000000000000000,
24'b000000010111000000010001,
24'b000000000000000000000000,
24'b000000011000000000010001,
24'b000000000000000000000000,
24'b000000011000000000010001,
24'b000000000000000000000000,
24'b000000011001000000010001,
24'b000000000000000000000000,
24'b000000011001000000010010,
24'b000000000000000000000000,
24'b000000011010000000010010,
24'b000000000000000000000000,
24'b000000011011000000010010,
24'b000000000000000000000000,
24'b000000011011000000010010,
24'b000000000000000000000000,
24'b000000011100000000010010,
24'b000000000000000000000000,
24'b000000011100000000010010,
24'b000000000000000000000000,
24'b000000011101000000010011,
24'b000000000000000000000000,
24'b000000011101000000010011,
24'b000000000000000000000000,
24'b000000011110000000010011,
24'b000000000000000000000000,
24'b000000011111000000010011,
24'b000000000000000000000000,
24'b000000100000000000010100,
24'b000000000000000000000000,
24'b000000100000000000010100,
24'b000000000000000000000000,
24'b000000100001000000010100,
24'b000000000000000000000000,
24'b000000100010000000010100,
24'b000000000000000000000000,
24'b000000100011000000010100,
24'b000000000000000000000000,
24'b000000100100000000010101,
24'b000000000000000000000000,
24'b000000100101000000010101,
24'b000000000000000000000000,
24'b000000100110000000010101,
24'b000000000000000000000000,
24'b000000100111000000010101,
24'b000000000000000000000000,
24'b000000101000000000010101,
24'b000000000000000000000000,
24'b000000101001000000010110,
24'b000000000000000000000000,
24'b000000101011000000010110,
24'b000000000000000000000000,
24'b000000101100000000010110,
24'b000000000000000000000000,
24'b000000101101000000010111,
24'b000000000000000000000000,
24'b000000101111000000010111,
24'b000000000000000000000000,
24'b000000110001000000010111,
24'b000000000000000000000000,
24'b000000110010000000011000,
24'b000000000000000000000000,
24'b000000110100000000011000,
24'b000000000000000000000000,
24'b000000110110000000011000,
24'b000000000000000000000000,
24'b000000111000000000011000,
24'b000000000000000000000000,
24'b000000111010000000011000,
24'b000000000000000000000000,
24'b000000111101000000011001,
24'b000000000000000000000000,
24'b000001000000000000011001,
24'b000000000000000000000000,
24'b000001000010000000011001,
24'b000000000000000000000000,
24'b000001000110000000011001,
24'b000000000000000000000000,
24'b000001001001000000011001,
24'b000000000000000000000000,
24'b000001001100000000011001,
24'b000000000000000000000000,
24'b000001010001000000011001,
24'b000000000000000000000000,
24'b000001010101000000011001,
24'b000000000000000000000000,
24'b000001011010000000011000,
24'b000000000000000000000000,
24'b000001100000000000010111,
24'b000000000000000000000000,
24'b000001100110000000010110,
24'b000000000000000000000000,
24'b000001101101000000010100,
24'b000000000000000000000000,
24'b000001110110000000010010,
24'b000000000000000000000000,
24'b000001111111000000001110,
24'b000000000000000000000000,
24'b000010001010000000001001,
24'b000000000000000000000000,
24'b000010010111000000000000,
24'b000000000000000000000000,
24'b000010100101111111110100,
24'b000000000000000000000000,
24'b000010110110111111011101,
24'b000000000000000000000000,
24'b000011000101111110110011,
24'b000000000000000000000000,
24'b000011000010111101001111,
24'b000000000000000000000000,
24'b111110110111110101110110,
24'b001111011111110000100001,
24'b011011010010000100000110,
24'b001111011111001111011111,
24'b001001001001010111000100,
24'b110000100001001111011111,
24'b000001001111110110000101,
24'b001111011111001111011111,
24'b110000110010010100011011,
24'b110000100001110000100001,
24'b010101100101110101011001,
24'b001111011111001111011111,
24'b000110000000010100101100,
24'b110000100001001111011110,
24'b000000110111110110100101,
24'b001111011111001111011111,
24'b111100101110010111110000,
24'b110000100001001111011111,
24'b110111011101000100101010,
24'b110000100001001111011111,
24'b100111100110110010001000,
24'b001111011111110000100001,
24'b001011101111010101110010,
24'b110000100001001111011111,
24'b111001011110000101000101,
24'b110000100001001111011111,
24'b100110001110111110000101,
24'b110000100001110000100001,
24'b000011010100110010101010,
24'b000000000000000000000000,
24'b000101101100111111111010,
24'b110000100001001111011111,
24'b110110001000100110100110,
24'b001111011111001111011111,
24'b100000100110111011001110,
24'b001111011111110000100001,
24'b110100010010000110000011,
24'b001111011111110000100001,
24'b111100001111011011100010,
24'b110000100001110000100001,
24'b000100000010001000010010,
24'b110000100001110000100001,
24'b010111001000000000111110,
24'b110000100001001111011111,
24'b000000000101111010001011,
24'b110000100010001111011111,
24'b101001011101101001010100,
24'b001111011111110000100001,
24'b111110101000001100100011,
24'b110000100001110000100001,
24'b010010111100111001001100,
24'b110000100010001111011111,
24'b110010101001100011111110,
24'b001111011111110000100001,
24'b010001111100111001000110,
24'b001111011111001111011111,
24'b111000010010001000010001,
24'b000000000000000000000000,
24'b111101101110000001011001,
24'b000000000000000000000000,
24'b111110100011000000001001,
24'b000000000000000000000000,
24'b111110110110111111101101,
24'b000000000000000000000000,
24'b111110111111111111100010,
24'b000000000000000000000000,
24'b111111000101111111011100,
24'b000000000000000000000000,
24'b111111001000111111011010,
24'b000000000000000000000000,
24'b111111001011111111011010,
24'b000000000000000000000000,
24'b111111001101111111011010,
24'b000000000000000000000000,
24'b111111001111111111011011,
24'b000000000000000000000000,
24'b111111010000111111011100,
24'b000000000000000000000000,
24'b111111010010111111011101,
24'b000000000000000000000000,
24'b111111010011111111011110,
24'b000000000000000000000000,
24'b111111010100111111011111,
24'b000000000000000000000000,
24'b111111010101111111100000,
24'b000000000000000000000000,
24'b111111010110111111100001,
24'b000000000000000000000000,
24'b111111010111111111100010,
24'b000000000000000000000000,
24'b111111011000111111100100,
24'b000000000000000000000000,
24'b111111011001111111100101,
24'b000000000000000000000000,
24'b111111011010111111100110,
24'b000000000000000000000000,
24'b111111011011111111100110,
24'b000000000000000000000000,
24'b111111011011111111100111,
24'b000000000000000000000000,
24'b111111011100111111101000,
24'b000000000000000000000000,
24'b111111011101111111101001,
24'b000000000000000000000000,
24'b111111011110111111101010,
24'b000000000000000000000000,
24'b111111011110111111101010,
24'b000000000000000000000000,
24'b111111011111111111101011,
24'b000000000000000000000000,
24'b111111011111111111101100,
24'b000000000000000000000000,
24'b111111100000111111101100,
24'b000000000000000000000000,
24'b111111100000111111101101,
24'b000000000000000000000000,
24'b111111100001111111101110,
24'b000000000000000000000000,
24'b111111100001111111101110,
24'b000000000000000000000000,
24'b111111100010111111101111,
24'b000000000000000000000000,
24'b111111100010111111101111,
24'b000000000000000000000000,
24'b111111100011111111101111,
24'b000000000000000000000000,
24'b111111100011111111110000,
24'b000000000000000000000000,
24'b111111100100111111110000,
24'b000000000000000000000000,
24'b111111100100111111110001,
24'b000000000000000000000000,
24'b111111100100111111110001,
24'b000000000000000000000000,
24'b111111100101111111110010,
24'b000000000000000000000000,
24'b111111100101111111110010,
24'b000000000000000000000000,
24'b111111100101111111110011,
24'b000000000000000000000000,
24'b111111100110111111110011,
24'b000000000000000000000000,
24'b111111100110111111110011,
24'b000000000000000000000000,
24'b111111100111111111110011,
24'b000000000000000000000000,
24'b111111100111111111110100,
24'b000000000000000000000000,
24'b111111100111111111110100,
24'b000000000000000000000000,
24'b111111101000111111110100,
24'b000000000000000000000000,
24'b111111101000111111110101,
24'b000000000000000000000000,
24'b111111101000111111110101,
24'b000000000000000000000000,
24'b111111101000111111110101,
24'b000000000000000000000000,
24'b111111101001111111110101,
24'b000000000000000000000000,
24'b111111101001111111110110,
24'b000000000000000000000000,
24'b111111101010111111110110,
24'b000000000000000000000000,
24'b111111101001111111110110,
24'b000000000000000000000000,
24'b111111101010111111110110,
24'b000000000000000000000000,
24'b111111101010111111110111,
24'b000000000000000000000000,
24'b111111101010111111110111,
24'b000000000000000000000000,
24'b111111101010111111110111,
24'b000000000000000000000000,
24'b111111101011111111110111,
24'b000000000000000000000000,
24'b111111101011111111110111,
24'b000000000000000000000000,
24'b111111101011111111111000,
24'b000000000000000000000000,
24'b111111101011111111111000,
24'b000000000000000000000000,
24'b111111101100111111111000,
24'b000000000000000000000000,
24'b111111101100111111111000,
24'b000000000000000000000000,
24'b111111101100111111111000,
24'b000000000000000000000000,
24'b111111101100111111111001,
24'b000000000000000000000000,
24'b111111101100111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111001,
24'b000000000000000000000000,
24'b111111101101111111111010,
24'b000000000000000000000000,
24'b111111101101111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101110111111111010,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111101111111111111011,
24'b000000000000000000000000,
24'b111111110000111111111011,
24'b000000000000000000000000,
24'b111111110000111111111011,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110000111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111100,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110001111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111101,
24'b000000000000000000000000,
24'b111111110010111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111101,
24'b000000000000000000000000,
24'b111111110011111111111101,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110011111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111110,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110100111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101111111111111,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110101000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110110000000000000,
24'b000000000000000000000000,
24'b111111110111000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000000,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111110111000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000001,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111000000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111001000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000010,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111010000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000011,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111011000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111100000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000100,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101,
24'b000000000000000000000000,
24'b111111111101000000000101};