logic pream_i [0:1559] = {
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
1,
0,
0,
1,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
0,
1,
0,
0,
0,
0,
1,
1,
1,
0,
0,
1,
0,
1,
0,
1,
0,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
1,
0,
1,
1,
0,
0,
1,
0,
1,
1,
0,
0,
1,
1,
1,
0,
0,
0,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
1,
1,
0,
0,
0,
0,
0,
0,
1,
1,
0,
0,
0,
0,
0,
0,
1,
1,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
0,
1,
0,
0,
1,
1,
1,
0,
0,
0,
1,
1,
0,
1,
1,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
0,
1,
1,
0,
0,
1,
1,
0,
1,
0,
0,
1,
1,
0,
1,
1,
0,
1,
1,
0,
1,
0,
0,
0,
1,
1,
0,
1,
1,
0,
0,
1,
1,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
1,
1,
0,
1,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
1,
0,
0,
0,
1,
1,
0,
0,
0,
0,
1,
1,
0,
1,
0,
1,
0,
1,
1,
0,
1,
1,
0,
0,
1,
0,
1,
1,
1,
0,
0,
1,
0,
1,
0,
0,
0,
1,
1,
1,
0,
1,
0,
1,
1,
0,
1,
0,
0,
1,
1,
1,
0,
1,
0,
1,
0,
1,
1,
1,
0,
0,
0,
1,
1,
1,
0,
1,
1,
1,
0,
0,
1,
0,
0,
1,
1,
0,
1,
1,
0,
1,
1,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
1,
1,
1,
0,
1,
0,
1,
0,
0,
0,
0,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
1,
0,
0,
0,
0,
0,
0,
1,
0,
1,
0,
0,
0,
0,
1,
0,
0,
0,
1,
1,
1,
1,
1,
1,
0,
1,
1,
1,
1,
0,
1,
0,
0,
1,
0,
1,
0,
1,
1,
0,
0,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
0,
1,
1,
0,
1,
0,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
1,
0,
0,
1,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
0,
1,
0,
0,
0,
0,
1,
1,
1,
0,
0,
1,
0,
1,
0,
1,
0,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
1,
0,
1,
1,
0,
0,
1,
0,
1,
1,
0,
0,
1,
1,
1,
0,
0,
0,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
1,
1,
0,
0,
0,
0,
0,
0,
1,
1,
0,
0,
0,
0,
0,
0,
1,
1,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
0,
1,
0,
0,
1,
1,
1,
0,
0,
0,
1,
1,
0,
1,
1,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
0,
1,
1,
0,
0,
1,
1,
0,
1,
0,
0,
1,
1,
0,
1,
1,
0,
1,
1,
0,
1,
0,
0,
0,
1,
1,
0,
1,
1,
0,
0,
1,
1,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
1,
1,
0,
1,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
1,
0,
0,
0,
1,
1,
0,
0,
0,
0,
1,
1,
0,
1,
0,
1,
0,
1,
1,
0,
1,
1,
0,
0,
1,
0,
1,
1,
1,
0,
0,
1,
0,
1,
0,
0,
0,
1,
1,
1,
0,
1,
0,
1,
1,
0,
1,
0,
0,
1,
1,
1,
0,
1,
0,
1,
0,
1,
1,
1,
0,
0,
0,
1,
1,
1,
0,
1,
1,
1,
0,
0,
1,
0,
0,
1,
1,
0,
1,
1,
0,
1,
1,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
1,
1,
1,
0,
1,
0,
1,
0,
0,
0,
0,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
1,
0,
0,
0,
0,
0,
0,
1,
0,
1,
0,
0,
0,
0,
1,
0,
0,
0,
1,
1,
1,
1,
1,
1,
0,
1,
1,
1,
1,
0,
1,
0,
0,
1,
0,
1,
0,
1,
1,
0,
0,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
0,
1,
1,
0,
1,
0,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
1,
0,
1,
1,
1,
0,
1,
0,
0,
1,
0,
0,
1,
0,
0,
0,
1,
1,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
1,
0,
0,
1,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
0,
1,
1,
1,
0,
1,
0,
0,
1,
0,
1,
0,
1,
1,
0,
1,
0,
0,
0,
1,
0,
0,
1,
0,
1,
1,
1,
1,
1,
0,
0,
0,
0,
0,
1,
0,
1,
1,
1,
1,
0,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
0,
1,
1,
0,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
1,
1,
0,
1,
0,
1,
1,
0,
0,
1,
1,
0,
0,
0,
1,
1,
1,
1,
0,
1,
0,
1,
1,
0,
0,
1,
1,
0,
0,
1,
1,
1,
0,
0,
0,
0,
1,
1,
1,
0,
0,
1,
0,
0,
1,
0,
0,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
1,
1,
1,
1,
1,
1,
0,
0,
1,
1,
1,
0,
1,
1,
1,
1,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
0,
0,
1,
0,
0,
1,
1,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
1,
1,
0,
1,
1,
1,
1,
0,
1,
1,
0,
1,
0,
1,
0,
0,
1,
1,
0,
0,
1,
0,
1,
1,
1,
1,
0,
0,
0,
0,
1,
0,
1,
1,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
0,
1,
0,
1,
1,
1,
0,
0,
1,
1,
0,
0,
0,
1,
1,
0,
1,
1,
1,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
1,
0,
1,
1,
1,
0,
0,
1,
1,
1,
1,
0,
1,
1,
1,
1,
0,
1,
0,
0,
0,
1,
1,
0,
1,
0,
1,
0,
1,
1,
1,
1,
1,
1,
0,
1,
0,
0,
1,
1,
0,
1,
1,
0,
0,
0,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
1,
1,
1,
1,
0,
1,
1,
0,
0,
0,
0,
1,
0,
1,
0,
1,
1,
0,
1,
1,
0,
0,
1,
0,
0,
1,
1,
1,
1,
1,
0,
1,
1,
1,
0,
1,
0,
0,
1,
0,
0,
1,
0,
0,
0,
1,
1,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
1,
0,
0,
1,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
0,
1,
1,
1,
0,
1,
0,
0,
1,
0,
1,
0,
1,
1,
0,
1,
0,
0,
0,
1,
0,
0,
1,
0,
1,
1,
1,
1,
1,
0,
0,
0,
0,
0,
1,
0,
1,
1,
1,
1,
0,
0,
0,
1,
1,
1,
1,
0,
0,
1,
1,
0,
1,
1,
0,
0,
1,
1,
1,
1,
1,
0,
1,
0,
1,
1,
1,
0,
1,
0,
1,
1,
0,
0,
1,
1,
0,
0,
0,
1,
1,
1,
1,
0,
1,
0,
1,
1,
0,
0,
1,
1,
0,
0,
1,
1,
1,
0,
0,
0,
0,
1,
1,
1,
0,
0,
1,
0,
0,
1,
0,
0,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
1,
1,
1,
1,
1,
1,
0,
0,
1,
1,
1,
0,
1,
1,
1,
1,
0,
0,
0,
0,
1,
1,
0,
0,
1,
0,
0,
0,
1,
0,
0,
1,
1,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
1,
1,
0,
1,
1,
1,
1,
0,
1,
1,
0,
1,
0,
1,
0,
0,
1,
1,
0,
0,
1,
0,
1,
1,
1,
1,
0,
0,
0,
0,
1,
0,
1,
1,
0,
0,
0,
1,
0,
1,
0,
1,
0,
1,
0,
1,
0,
1,
1,
1,
0,
0,
1,
1,
0,
0,
0,
1,
1,
0,
1,
1,
1,
0,
1,
1,
1,
0,
1,
1,
1,
1,
1,
1,
0,
1,
1,
1,
0,
0,
1,
1,
1,
1,
0,
1,
1,
1,
1,
0,
1,
0,
0,
0,
1,
1,
0,
1,
0,
1,
0,
1,
1,
1,
1,
1,
1,
0,
1,
0,
0,
1,
1,
0,
1,
1,
0,
0,
0,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
1,
1,
1,
1,
0,
1,
1,
0,
0,
0,
0,
1,
0,
1,
0,
1,
1,
0,
1,
1,
0,
0,
1,
0,
0,
1,
1,
1};