logic [13:0] addr_rand_interl [0:4607] = {
14'b00111111001001,
14'b00100110101010,
14'b00100101111110,
14'b00100111101111,
14'b00000011011011,
14'b00100010101110,
14'b00001001000111,
14'b00101101100001,
14'b00000100111100,
14'b00111101000100,
14'b00110101101111,
14'b00100011011000,
14'b00011011110010,
14'b01000010011001,
14'b00000011110101,
14'b00001010011000,
14'b01000001110000,
14'b01000001011000,
14'b00010100000100,
14'b00011110101101,
14'b00101100101010,
14'b00011001010110,
14'b00000101100110,
14'b00001000101100,
14'b00101111100001,
14'b00100010100101,
14'b00011000010101,
14'b00010000010111,
14'b00110000010100,
14'b00001101011101,
14'b00110110010110,
14'b00111000110010,
14'b00100110010010,
14'b01000010010110,
14'b00111111111001,
14'b00111110110101,
14'b00010010110000,
14'b00100101011111,
14'b00110100100010,
14'b00000101111111,
14'b00001011000110,
14'b00011011011000,
14'b00100111100011,
14'b01000101110101,
14'b00111101001101,
14'b00000110111111,
14'b00000111101001,
14'b00110101101001,
14'b00010111101100,
14'b00010010011110,
14'b00011111000000,
14'b00110111101001,
14'b00100111001110,
14'b00101011110011,
14'b00100010110110,
14'b00111010011110,
14'b00100001000110,
14'b00110001101101,
14'b00001001010100,
14'b00100100010000,
14'b00000111111111,
14'b00100010100000,
14'b00001100011001,
14'b00110011110100,
14'b00100010011011,
14'b00001011000100,
14'b00010001001110,
14'b00100000111011,
14'b00001011000010,
14'b01000000101101,
14'b00101000010001,
14'b00100110101101,
14'b01000100001110,
14'b00010111110000,
14'b00110000110100,
14'b00010010111000,
14'b00001100001110,
14'b00001000010010,
14'b00011000011100,
14'b00100000100110,
14'b00011000110010,
14'b00000101110011,
14'b00001101010101,
14'b00010010010001,
14'b00101001111011,
14'b00010110101011,
14'b00111010110011,
14'b00100111010001,
14'b00101000010101,
14'b00110010010110,
14'b00100101100010,
14'b00000000010001,
14'b00111010000111,
14'b00011011111000,
14'b00011111001101,
14'b00010011101101,
14'b00111011010110,
14'b01000001101101,
14'b00110110100100,
14'b00011011111100,
14'b00010100001011,
14'b00100101011000,
14'b00101101101100,
14'b00101101000101,
14'b00101100011001,
14'b00101100110100,
14'b01000001000100,
14'b00000110101001,
14'b00110101111010,
14'b00101010110100,
14'b00000000001011,
14'b00000011011100,
14'b01000110111010,
14'b00001011100110,
14'b00101100011011,
14'b00011101010000,
14'b00111010000011,
14'b00101011000110,
14'b00010010010010,
14'b00101101001100,
14'b00010011100101,
14'b00011000111110,
14'b00100011001101,
14'b00011001011010,
14'b00110011101101,
14'b00010011110000,
14'b00110000101100,
14'b00001111100111,
14'b00100010011010,
14'b00101010011000,
14'b00111111110011,
14'b00111100110001,
14'b00100000111100,
14'b00110111100100,
14'b00110100111001,
14'b00101101011000,
14'b00111011101111,
14'b00101010000011,
14'b00110101001000,
14'b00110101010101,
14'b00001010101010,
14'b00110010110010,
14'b00111111011110,
14'b00110100000011,
14'b01000001010011,
14'b01000011101111,
14'b00001100000011,
14'b00111101011001,
14'b01000101000010,
14'b00100011000000,
14'b00110111011111,
14'b00010100011001,
14'b00110110000101,
14'b00000101010001,
14'b01000011110000,
14'b00100101011010,
14'b00011011000001,
14'b01000110001110,
14'b00011011001001,
14'b00010011100010,
14'b00101011011101,
14'b00011011000100,
14'b00000101011111,
14'b00011000010111,
14'b00101110001011,
14'b00000011110011,
14'b00000100000011,
14'b00111011100101,
14'b00011000110001,
14'b00101001110001,
14'b00100011100000,
14'b00011111101110,
14'b00110011000010,
14'b01000110100100,
14'b00110000110110,
14'b00011010000100,
14'b00001001011000,
14'b00011100011100,
14'b00001011110101,
14'b01000011011101,
14'b00010100110110,
14'b00011001011011,
14'b00000010111011,
14'b01000011011001,
14'b00101110000111,
14'b01000100110100,
14'b00000011100100,
14'b00110111101100,
14'b00101110010111,
14'b00010110010101,
14'b00100001101101,
14'b00110011110111,
14'b00100010011111,
14'b00110010110000,
14'b00100111100100,
14'b00100001001001,
14'b00011000011101,
14'b00000101001110,
14'b00000001111000,
14'b01000010001100,
14'b01000100110110,
14'b00001010111110,
14'b00001010101110,
14'b00100110011101,
14'b01000011001111,
14'b01000111100101,
14'b01000011011010,
14'b00000101011001,
14'b00011110100101,
14'b00000000001001,
14'b00011001010100,
14'b00001100010010,
14'b00100100111011,
14'b00010001011001,
14'b00011000001110,
14'b00100101100100,
14'b00011101011000,
14'b00001110100000,
14'b00110101000111,
14'b00001101011110,
14'b00101000011101,
14'b00000010111100,
14'b00000111111101,
14'b00110001001111,
14'b00000100010010,
14'b00000010000010,
14'b00110101111101,
14'b00101000010000,
14'b00110010101011,
14'b00101011001110,
14'b00100101101101,
14'b00111110010011,
14'b00010000110010,
14'b00110011100100,
14'b00110101001110,
14'b01000110011110,
14'b00100101111100,
14'b00110101011110,
14'b00001111010100,
14'b00010100100000,
14'b00011110001111,
14'b01000101101010,
14'b00110100101001,
14'b00000110101101,
14'b00010111100101,
14'b00011010111110,
14'b00000001000011,
14'b00000011111000,
14'b00110110101001,
14'b01000110010100,
14'b00000011000110,
14'b00100100011000,
14'b01000111111100,
14'b00111001100111,
14'b00110110110111,
14'b00100110110110,
14'b00110100101111,
14'b01000000011101,
14'b00010101100000,
14'b00000010001100,
14'b00011110001110,
14'b00010110111001,
14'b00100000000111,
14'b00011100000010,
14'b00111100011011,
14'b00101110101110,
14'b00001010111001,
14'b00010010001111,
14'b00100111101100,
14'b00011100101000,
14'b00100000110010,
14'b00001000000111,
14'b00111001111111,
14'b01000101011100,
14'b00000001001100,
14'b00001100101011,
14'b00111011001000,
14'b00011000001100,
14'b00110000011101,
14'b00010110101111,
14'b00100110100010,
14'b00011110001010,
14'b00110100000101,
14'b00000011001001,
14'b00010100010111,
14'b01000100000100,
14'b00010100011000,
14'b00101101110001,
14'b00000111001001,
14'b00000010000001,
14'b00101100001000,
14'b00111001101001,
14'b00100101111010,
14'b00100000101100,
14'b00110111000000,
14'b00111110111101,
14'b00100011001000,
14'b01000100110010,
14'b00011011101001,
14'b00101011100011,
14'b01000100110111,
14'b00000001001101,
14'b00010111000000,
14'b00000100101000,
14'b00011001110010,
14'b00101001001110,
14'b01000100001011,
14'b00011111111110,
14'b00000001110011,
14'b00010011101010,
14'b00011111100110,
14'b00110110110010,
14'b00000011000100,
14'b01000101010110,
14'b00011011111110,
14'b00100011100111,
14'b01000101011110,
14'b00111101010011,
14'b00010010010100,
14'b00001111111010,
14'b00000011001100,
14'b00101110001101,
14'b00100010101000,
14'b00110111111110,
14'b00000011001010,
14'b00010111011111,
14'b00110111001011,
14'b00011011010000,
14'b00100100011010,
14'b00010001001100,
14'b00111000001011,
14'b00101010000010,
14'b00001010011111,
14'b00100010111000,
14'b00111110010001,
14'b00101001101101,
14'b00100101101000,
14'b00001011010101,
14'b00001000111111,
14'b00100011111000,
14'b00101011100111,
14'b00010010000101,
14'b00100010000000,
14'b00011010001110,
14'b00011010011101,
14'b00110110001001,
14'b00111101010110,
14'b00001100100100,
14'b00000111110011,
14'b00001010100100,
14'b01000100000110,
14'b01000101101101,
14'b00100111010100,
14'b00100110101001,
14'b00101000001000,
14'b00111010101101,
14'b01000100010111,
14'b00111101111110,
14'b00000110100011,
14'b00101000110110,
14'b00111111000011,
14'b00001111111000,
14'b01000000000010,
14'b00100001001011,
14'b00110010011101,
14'b00000010000011,
14'b01000010101011,
14'b00110010110001,
14'b00110011001101,
14'b00101111011011,
14'b00100011101100,
14'b00000100101110,
14'b00000110001010,
14'b00100110010011,
14'b00010000001101,
14'b00111011110111,
14'b00001011010100,
14'b00010110001111,
14'b00111010110110,
14'b00001001001001,
14'b00010110000100,
14'b00011111110100,
14'b00101001011001,
14'b00000111010010,
14'b00011011000101,
14'b00000000110110,
14'b00111100100010,
14'b00101110000100,
14'b01000100000001,
14'b00101101010011,
14'b00100111010111,
14'b00111001110110,
14'b00101001010000,
14'b00011101110101,
14'b00000100111000,
14'b00011000010100,
14'b00000001101011,
14'b00101011101100,
14'b00010110000110,
14'b00111001101010,
14'b00111100000001,
14'b00010111010011,
14'b00100001100100,
14'b00101011000111,
14'b00101010100000,
14'b00100110101110,
14'b00000010101000,
14'b00000000100100,
14'b01000001110100,
14'b00110100000000,
14'b00100000010010,
14'b00001001010000,
14'b00001000110100,
14'b00101100111100,
14'b00001110011010,
14'b00101101110100,
14'b00001101001111,
14'b00110011001000,
14'b00010101011100,
14'b00101101100110,
14'b01000001100110,
14'b00000010110000,
14'b00111000100111,
14'b00100101100111,
14'b00011100011011,
14'b00100001101110,
14'b00011100000100,
14'b01000101001100,
14'b00001110101100,
14'b00111100111000,
14'b00111001011100,
14'b00111001010110,
14'b00010100010010,
14'b00001001110101,
14'b00011010101100,
14'b00100111010000,
14'b00101100101011,
14'b01000011110111,
14'b01000001010111,
14'b00101101101000,
14'b00010001000011,
14'b00000001010000,
14'b00001010000011,
14'b00011001101111,
14'b00101011010011,
14'b00101101010000,
14'b00000100111010,
14'b00101111110101,
14'b00010010110100,
14'b00110000011110,
14'b00011110101111,
14'b00110100010110,
14'b00001100011000,
14'b00100100011111,
14'b00101100101111,
14'b00111101110110,
14'b00010010011010,
14'b00101010111000,
14'b01000001111101,
14'b00111100011001,
14'b00101010011111,
14'b00000111110101,
14'b00111000110011,
14'b00101001000011,
14'b00000111001100,
14'b01000000011110,
14'b00101000111100,
14'b00010110100111,
14'b00011111011110,
14'b00111101010111,
14'b00000111000110,
14'b00001111001100,
14'b00001101010000,
14'b00001011111111,
14'b00101100110101,
14'b00101110100001,
14'b00101111110100,
14'b00100110110101,
14'b00010001111110,
14'b00100001011101,
14'b01000010101001,
14'b00100001011001,
14'b00101100111011,
14'b00011001000001,
14'b00010010001011,
14'b00101111001010,
14'b00011011101111,
14'b00111101000101,
14'b00101100000011,
14'b00111001000111,
14'b01000000001111,
14'b01000110010110,
14'b00111101100110,
14'b00000100001010,
14'b01000000001001,
14'b01000111110000,
14'b01000101001110,
14'b00101011110010,
14'b00000100100011,
14'b00110001100010,
14'b00101110111001,
14'b00010011010111,
14'b00101100111111,
14'b00001111011010,
14'b01000111111000,
14'b00101110000110,
14'b01000010001010,
14'b00111011010100,
14'b00001001111101,
14'b00010011001000,
14'b00010101101001,
14'b00101100010101,
14'b00100011110001,
14'b00101100000101,
14'b00001000001001,
14'b01000100010100,
14'b00110101101010,
14'b00010110001101,
14'b01000010011110,
14'b00111110100111,
14'b00011101100100,
14'b00010100010110,
14'b00000101100000,
14'b00100100001111,
14'b01000011000111,
14'b01000001110001,
14'b01000100110101,
14'b00011011110110,
14'b00100010000101,
14'b00101110010011,
14'b00001111100011,
14'b00101100000010,
14'b00101001010110,
14'b00110000000010,
14'b00010101010111,
14'b00010001111001,
14'b00100110000001,
14'b00110101000001,
14'b00101110111110,
14'b00101111101100,
14'b00011100010101,
14'b00010000100011,
14'b00100111011100,
14'b00010001011011,
14'b00011010111001,
14'b00011000111101,
14'b00111111000101,
14'b00111101100101,
14'b00011001111110,
14'b00001111101000,
14'b00001001111001,
14'b00011010110111,
14'b00001010000101,
14'b00000000000111,
14'b00110100011000,
14'b00111100001000,
14'b00000100100111,
14'b00100000000000,
14'b00011001100011,
14'b01000011010010,
14'b00010011111100,
14'b00100011000010,
14'b00110100100110,
14'b00001000101000,
14'b00111101111000,
14'b00000111100000,
14'b00100110001011,
14'b00110110101100,
14'b00010111001001,
14'b00101101001111,
14'b00000001010001,
14'b00100001010100,
14'b01000110111101,
14'b00011110111111,
14'b00010110001010,
14'b00110001100011,
14'b00010011100000,
14'b00011000111000,
14'b00110011010101,
14'b00100001110101,
14'b00010001000111,
14'b00010101110101,
14'b00010011001010,
14'b00110000000000,
14'b00001101011010,
14'b00010101111010,
14'b01000011111011,
14'b00000011101000,
14'b00001001000101,
14'b01000100010110,
14'b00111101110101,
14'b00011111111000,
14'b00101010010110,
14'b00011111101001,
14'b00010101010001,
14'b00110010110111,
14'b00111111001100,
14'b00111010001010,
14'b01000010010010,
14'b00000100111011,
14'b00100100100101,
14'b00111011001101,
14'b00011001101000,
14'b00000101011110,
14'b00100111000011,
14'b00100011000110,
14'b00101111000010,
14'b00111111010011,
14'b00000010010110,
14'b00011111011100,
14'b00010001011010,
14'b01000111100100,
14'b00100001001100,
14'b01000100111000,
14'b00011101010111,
14'b01000101000111,
14'b00001011111001,
14'b00111101011010,
14'b01000001001000,
14'b00111101111001,
14'b00010110000111,
14'b01000111001000,
14'b00111100110101,
14'b00111111010111,
14'b00101000000110,
14'b00000110111010,
14'b00111001011101,
14'b00101010001011,
14'b00010101001000,
14'b00100000111001,
14'b00101101000110,
14'b00001000111101,
14'b00001000100100,
14'b00011011111001,
14'b00000001110110,
14'b00110111011010,
14'b00011010000001,
14'b00110110000011,
14'b00010000100101,
14'b00011011111010,
14'b00011101110111,
14'b00110000111011,
14'b00110000100110,
14'b00000110100101,
14'b00000011101111,
14'b00000101001011,
14'b00101010100010,
14'b00010000011001,
14'b00001001111010,
14'b00101100111110,
14'b01000111000101,
14'b00001011011100,
14'b00010101110010,
14'b00111000011111,
14'b00011001110001,
14'b00111010010001,
14'b00101001110101,
14'b00010111001100,
14'b00001000010000,
14'b00010011000001,
14'b00111000111001,
14'b00110111100101,
14'b00110100001110,
14'b00100110111000,
14'b00010111100100,
14'b00110100001001,
14'b00000001001111,
14'b00010100000101,
14'b00100000010100,
14'b01000000111001,
14'b00000101111101,
14'b00100010101010,
14'b00101100010010,
14'b00000011010111,
14'b00101111111100,
14'b00110111101110,
14'b01000010101101,
14'b00011100110110,
14'b00000010011010,
14'b00101001010101,
14'b00100001100101,
14'b01000011011110,
14'b00101111101010,
14'b00100000110011,
14'b00101011101101,
14'b00111000100110,
14'b00011111101000,
14'b00011011100111,
14'b00101010100001,
14'b00001010011011,
14'b00001100010110,
14'b00000011000000,
14'b00101000010111,
14'b01000111000111,
14'b00000000011000,
14'b01000000010011,
14'b01000101111110,
14'b00000110101000,
14'b00000011010100,
14'b01000111011000,
14'b00001000000010,
14'b00100100110011,
14'b01000100101100,
14'b00000010010000,
14'b00111010000110,
14'b01000011100111,
14'b00001000001000,
14'b00110001101010,
14'b00110011011111,
14'b01000011000001,
14'b00100010001010,
14'b01000101110100,
14'b00111111101010,
14'b00101101101111,
14'b00110010100111,
14'b00110101001010,
14'b00111111001011,
14'b00111001001011,
14'b00001011110001,
14'b00100100111111,
14'b00011100001111,
14'b00100100101011,
14'b00010110100001,
14'b00001010001011,
14'b00101101111010,
14'b01000101101110,
14'b00000011011110,
14'b00101010101010,
14'b00111101111100,
14'b01000111011100,
14'b00110111000001,
14'b01000011111000,
14'b00000111101000,
14'b00001100001011,
14'b00110110111100,
14'b01000010111101,
14'b00001011011101,
14'b00110011010100,
14'b00111101000010,
14'b00111111101100,
14'b00001110101001,
14'b00100101001011,
14'b00100010001101,
14'b01000100100010,
14'b00100110101000,
14'b00010101100010,
14'b00011001101011,
14'b00100011100110,
14'b00001101111101,
14'b00111011011101,
14'b01000111011011,
14'b00011101010101,
14'b00101101000011,
14'b00000101110101,
14'b00010110001100,
14'b00000010000111,
14'b00011100000111,
14'b00101010101100,
14'b00101010001101,
14'b00100110110001,
14'b00011001100010,
14'b00110100011110,
14'b00111101011110,
14'b00010111111011,
14'b00110000010111,
14'b00011001010000,
14'b00001110010100,
14'b00000100000001,
14'b00000111001111,
14'b00100000100111,
14'b00100001000010,
14'b00001011000101,
14'b00000100100101,
14'b01000010000001,
14'b00001101000010,
14'b01000000110010,
14'b00110001110010,
14'b00010100111111,
14'b00110000111001,
14'b00111100010110,
14'b00000111001101,
14'b01000111101101,
14'b00010111110001,
14'b00001110111110,
14'b00111011110011,
14'b00000111100110,
14'b00001000000101,
14'b01000011010011,
14'b00011001000111,
14'b00111100110011,
14'b01000110110001,
14'b00101110001000,
14'b00011101111111,
14'b00111101000001,
14'b00000001110010,
14'b00010100111110,
14'b00011111010101,
14'b00011000010011,
14'b00010110000001,
14'b00110101010001,
14'b00000110101110,
14'b00010001110110,
14'b00100101100000,
14'b00101000001010,
14'b00111101011011,
14'b00101100111000,
14'b00111110001011,
14'b00100110000110,
14'b00001001001010,
14'b00111100101000,
14'b00100101110010,
14'b01000011110100,
14'b01000100100001,
14'b00111100100011,
14'b01000100000101,
14'b00010111011011,
14'b00100001011000,
14'b01000111110011,
14'b01000100101001,
14'b00110111010101,
14'b00010001100001,
14'b01000000111111,
14'b01000010100000,
14'b00101100000100,
14'b00010111001101,
14'b00100011111001,
14'b00000011001101,
14'b00001010010100,
14'b01000101001010,
14'b00001110010101,
14'b00101101110000,
14'b00100101001101,
14'b00111001110010,
14'b00001001100100,
14'b00001101101111,
14'b00111001100010,
14'b00011011101000,
14'b00100001000000,
14'b00101010001100,
14'b00110010001011,
14'b00001010111101,
14'b01000100111111,
14'b00101110011110,
14'b00010100101001,
14'b00110001101011,
14'b00000001010011,
14'b00101101000010,
14'b00110000011011,
14'b00011101000000,
14'b00011001110101,
14'b00101100010001,
14'b00111101111101,
14'b01000110000000,
14'b00001111111100,
14'b00010100111101,
14'b00111110000111,
14'b00100010101011,
14'b01000111101110,
14'b00011101100101,
14'b01000010010001,
14'b00100001010111,
14'b00100011101110,
14'b00111001110000,
14'b00011010011011,
14'b00101000111110,
14'b00110110010101,
14'b00010101011000,
14'b01000110101000,
14'b00001111001111,
14'b00000001100101,
14'b00110100011010,
14'b00100011001011,
14'b00010110110001,
14'b00000101100001,
14'b00111101001111,
14'b00100010111011,
14'b00101110111000,
14'b00110011000110,
14'b00100100010010,
14'b01000111100010,
14'b00010100000110,
14'b00001100100010,
14'b00010101000111,
14'b01000100101110,
14'b00001011010000,
14'b00100000101101,
14'b00011110011100,
14'b00010111001110,
14'b00101111100100,
14'b00011111001011,
14'b00101110110111,
14'b00100010010111,
14'b00111000110111,
14'b00010010111101,
14'b00000001100100,
14'b00000101101011,
14'b00101101011111,
14'b00100001100111,
14'b00110101011100,
14'b00101010101001,
14'b01000010000011,
14'b00001101101011,
14'b00110110001101,
14'b00101011011011,
14'b00010010101100,
14'b01000001101111,
14'b00010101001110,
14'b00000001001110,
14'b00110111101000,
14'b00101000111010,
14'b01000011100101,
14'b00110011101110,
14'b00001111000010,
14'b00100000111101,
14'b00100000110111,
14'b00000000110100,
14'b00010100111010,
14'b00101011110110,
14'b00101100101101,
14'b00100011011011,
14'b00011010010011,
14'b00101001000001,
14'b00011010001100,
14'b00110001101000,
14'b00000101101111,
14'b00010000100100,
14'b00001011100011,
14'b00100110100000,
14'b00111000101000,
14'b00101000110111,
14'b00110111000010,
14'b00111001001111,
14'b00000010011111,
14'b00101000100110,
14'b00000000110011,
14'b01000101110011,
14'b00011111100101,
14'b00111111011001,
14'b00111111100101,
14'b00110001110011,
14'b00011000101010,
14'b00001001010010,
14'b01000111100001,
14'b00011100010010,
14'b00000000001000,
14'b00100001010001,
14'b01000010111000,
14'b00110000110011,
14'b00001111001001,
14'b01000010110100,
14'b00010001011100,
14'b00011011111101,
14'b00010111111000,
14'b00011100111000,
14'b00011111001110,
14'b00000001111001,
14'b00110111111100,
14'b00000110001111,
14'b00110110000000,
14'b00000100111101,
14'b00100111111010,
14'b00101101111001,
14'b00001101101110,
14'b01000100111011,
14'b00110111010000,
14'b00111001110011,
14'b00011111110101,
14'b00011111110001,
14'b00110111100001,
14'b00111011111100,
14'b00100100111100,
14'b00110001110001,
14'b00000111011001,
14'b00111001000000,
14'b00001001101110,
14'b00110101000000,
14'b00010001110010,
14'b00100110010110,
14'b00101000100010,
14'b01000101011111,
14'b00101101111101,
14'b00001110101000,
14'b00101110011010,
14'b00000010101001,
14'b00010110111101,
14'b00100101111001,
14'b00101000001011,
14'b00100110010100,
14'b01000101100110,
14'b00101010100100,
14'b00110000100010,
14'b00101000011011,
14'b00000100111110,
14'b00011011100010,
14'b00110001011100,
14'b00111001111011,
14'b00101110110011,
14'b00010110000000,
14'b00100100110000,
14'b01000011100000,
14'b00011010000011,
14'b00011001101100,
14'b00000001110001,
14'b00111101001001,
14'b00001101110100,
14'b00111000010111,
14'b00011110100111,
14'b00101100101100,
14'b00111100001101,
14'b00100110000111,
14'b00110001100101,
14'b00010111000110,
14'b00110010011010,
14'b01000101001011,
14'b00001000100110,
14'b00000100001110,
14'b00001011011001,
14'b00011101110011,
14'b00101100101110,
14'b01000011011011,
14'b01000001011110,
14'b01000110011011,
14'b00000000011100,
14'b01000000100001,
14'b01000011010111,
14'b00111100100111,
14'b00001110001111,
14'b00010011011101,
14'b00011001111100,
14'b00000011011000,
14'b00111100100001,
14'b00100001000001,
14'b00101111100010,
14'b00100010010101,
14'b00011010111010,
14'b00001101101100,
14'b00010101110001,
14'b00100110100111,
14'b00000000101000,
14'b00100010000111,
14'b00010000111000,
14'b00010010100111,
14'b01000110000010,
14'b00111010100001,
14'b00110010100011,
14'b00110101011010,
14'b00011110101110,
14'b00110100101011,
14'b00000011101001,
14'b00110000111010,
14'b00110111001000,
14'b01000011111111,
14'b00010111010110,
14'b00010110010010,
14'b00110010111010,
14'b00101011000010,
14'b00000001000110,
14'b00011110100000,
14'b00000010110100,
14'b00011000010010,
14'b00101101111000,
14'b00010000101000,
14'b00010000110011,
14'b00101011100100,
14'b00101001111001,
14'b00011100000011,
14'b00101001010011,
14'b00001110000111,
14'b00101001110000,
14'b00010011111111,
14'b00100111111111,
14'b00011010100100,
14'b00011100100101,
14'b01000010101000,
14'b01000000010111,
14'b00001110111010,
14'b00100010010110,
14'b00011000101110,
14'b00000111100111,
14'b00111100010101,
14'b00100001110011,
14'b00010111000010,
14'b00100100100111,
14'b00101000000111,
14'b00010111000111,
14'b00010001000010,
14'b00001001011010,
14'b00001111100010,
14'b00001010000010,
14'b00100101111011,
14'b00101110000001,
14'b00111000111100,
14'b00110011010111,
14'b00110110011110,
14'b00100011111110,
14'b00100101101100,
14'b00100001010101,
14'b01000111011110,
14'b00101100011010,
14'b00110110110110,
14'b00001111100100,
14'b00000010100000,
14'b00101110010101,
14'b00110000011111,
14'b00100010100010,
14'b00101100011000,
14'b00111000100100,
14'b00101000000010,
14'b00100000011100,
14'b00011110011101,
14'b00111010101000,
14'b00000001000100,
14'b00000011011001,
14'b00011101011101,
14'b00100001011110,
14'b00110100110001,
14'b00111000110001,
14'b01000100101010,
14'b00110101111110,
14'b00101001100100,
14'b00111001101101,
14'b00100010101100,
14'b00100001001000,
14'b00101011110100,
14'b00001001001011,
14'b00110111001001,
14'b00001000000110,
14'b00001000111010,
14'b00110000010011,
14'b00100001100000,
14'b00111110011010,
14'b00011001100100,
14'b00011000111111,
14'b00110100011111,
14'b00000011110110,
14'b00111101101111,
14'b00110011000101,
14'b00010111100001,
14'b00001110000001,
14'b00011110101100,
14'b01000001011111,
14'b00100111010101,
14'b00110101111100,
14'b00101011100010,
14'b00110000100011,
14'b01000100000000,
14'b00010111111101,
14'b00010101111011,
14'b00101100000111,
14'b00001100101110,
14'b00001000101110,
14'b00111100011110,
14'b00111111110111,
14'b01000110011101,
14'b00001011101101,
14'b00100011010010,
14'b00000100011110,
14'b00101101001000,
14'b00100011011100,
14'b00010011000101,
14'b00101111100000,
14'b00001001011001,
14'b00011101000101,
14'b00010011111110,
14'b00000100001111,
14'b00010111011101,
14'b00010011001001,
14'b00100101111000,
14'b00011000001001,
14'b00011111100010,
14'b00011100001001,
14'b00010100010101,
14'b00110011011010,
14'b01000110011001,
14'b00001111111001,
14'b00110101101101,
14'b00110010000011,
14'b01000100010101,
14'b01000001010001,
14'b00101111100111,
14'b00111000101011,
14'b00011110110110,
14'b00111000100101,
14'b01000111110001,
14'b00110100010001,
14'b00101100001101,
14'b00001100111110,
14'b01000111110100,
14'b00110100001101,
14'b00111001001010,
14'b00011000000100,
14'b00111111101101,
14'b00011010101111,
14'b00110110000010,
14'b00111010001101,
14'b00111110011111,
14'b00000000010011,
14'b00001001100110,
14'b00110010111101,
14'b00100000111010,
14'b00111010011101,
14'b00000010001000,
14'b00101000000011,
14'b00100101110110,
14'b00110100100001,
14'b00010000110111,
14'b00001110110001,
14'b00001000111000,
14'b00001110111111,
14'b00110110010111,
14'b00010110100100,
14'b01000110101001,
14'b00010111001011,
14'b01000010111111,
14'b00011110011111,
14'b00001001011100,
14'b00111101100010,
14'b00010000111010,
14'b00000001011000,
14'b00011110111011,
14'b00000011101011,
14'b00100111001011,
14'b00001111011011,
14'b00010010111010,
14'b00111000101010,
14'b00001001000110,
14'b00001100111100,
14'b00010010111111,
14'b00001001011011,
14'b00010000100111,
14'b00110111010010,
14'b00101010011100,
14'b00000000101011,
14'b00110101101000,
14'b00011011010100,
14'b01000011100110,
14'b00100001111000,
14'b00011111111001,
14'b00111011000011,
14'b00110101001011,
14'b00101111100101,
14'b00110001111110,
14'b00000101001000,
14'b00011100111011,
14'b00100011011101,
14'b00110011110000,
14'b00111101101000,
14'b00101001011000,
14'b01000000110011,
14'b00011110101000,
14'b00011111101101,
14'b00110001000101,
14'b00010101101100,
14'b00001111001000,
14'b00001000010111,
14'b00000001111101,
14'b00100111000101,
14'b00110110111000,
14'b00011111111010,
14'b00000011010101,
14'b00000011101110,
14'b00010100100010,
14'b01000100011001,
14'b00111010001100,
14'b00100011110000,
14'b00100111101000,
14'b00101111101111,
14'b01000011111100,
14'b00111100110000,
14'b00110110001010,
14'b00111111101111,
14'b00001011111100,
14'b00101111000111,
14'b00110010010010,
14'b00000000110001,
14'b00000000001110,
14'b00001110110110,
14'b00110000000111,
14'b00110010000111,
14'b00011001100110,
14'b00101100010011,
14'b00000010101101,
14'b00001010101101,
14'b00111000011001,
14'b00100101001001,
14'b00101001011011,
14'b00110101100011,
14'b00110101001001,
14'b00010011101000,
14'b01000100100000,
14'b00010100001111,
14'b00111011101000,
14'b00001010001000,
14'b00001111101001,
14'b00001111010011,
14'b00111101001011,
14'b00111010101001,
14'b00101000101001,
14'b00111011010010,
14'b00010111111001,
14'b00111110011110,
14'b01000000000011,
14'b00010001000001,
14'b00010101000110,
14'b01000010001111,
14'b01000000101010,
14'b00110110001100,
14'b00011000011000,
14'b00111100101100,
14'b00011111101010,
14'b00100101010110,
14'b00110011110001,
14'b00011011111011,
14'b00000000110000,
14'b00000000010101,
14'b00000110001101,
14'b00100101101001,
14'b00001000011110,
14'b00111100011100,
14'b00110100010101,
14'b00100011110110,
14'b00010110111100,
14'b00100001110001,
14'b01000011011000,
14'b00101010000001,
14'b00110100110011,
14'b00111010110101,
14'b00111011010001,
14'b00110000111000,
14'b00111001011110,
14'b00100110001100,
14'b00001110010111,
14'b00111111010001,
14'b00000010100101,
14'b00001110110010,
14'b00001101110000,
14'b00011000101100,
14'b00001010101100,
14'b00011001011111,
14'b01000101011010,
14'b00001100111010,
14'b00111111100100,
14'b00010010001000,
14'b00010100100100,
14'b00101101010101,
14'b00001100110001,
14'b00100001011111,
14'b00011110110100,
14'b00001001101001,
14'b00001110111000,
14'b00011110111001,
14'b00000100011001,
14'b00001000001010,
14'b00000010001110,
14'b00000000000011,
14'b00000110100100,
14'b00010010000000,
14'b00001010110101,
14'b00110111010111,
14'b00100111001001,
14'b00000000101100,
14'b00000101111001,
14'b00000101111010,
14'b00101110001110,
14'b00000110000001,
14'b00111101001000,
14'b00111000101100,
14'b00111000010101,
14'b00101111111001,
14'b01000101100111,
14'b00001010010010,
14'b00010011001011,
14'b00100000110001,
14'b00001101001000,
14'b00011001101110,
14'b00011010100111,
14'b00000011111001,
14'b00001010110110,
14'b00001011100001,
14'b00010100110010,
14'b00100110110111,
14'b00100110111100,
14'b00000111100010,
14'b00100111110111,
14'b00001100101010,
14'b00001000010110,
14'b00100011101010,
14'b01000000001101,
14'b00101010110010,
14'b00001111010110,
14'b00111010101110,
14'b00111010110111,
14'b00001100011101,
14'b00110011100110,
14'b00011110000101,
14'b01000001001110,
14'b00101011110111,
14'b00010110011001,
14'b00100101100011,
14'b01000111001011,
14'b00100111000001,
14'b00100011111111,
14'b00101111101000,
14'b00110010111001,
14'b00010101111111,
14'b00010000101010,
14'b00101100010000,
14'b00111011010111,
14'b00011000110011,
14'b00101001100011,
14'b00111111010101,
14'b00110101000110,
14'b00011010110101,
14'b00111110001100,
14'b00010110011011,
14'b00000101001111,
14'b00100000010111,
14'b00110000010000,
14'b00001100100001,
14'b00100111000000,
14'b00010000100000,
14'b00110101010111,
14'b00001011101011,
14'b01000000001011,
14'b00011001111101,
14'b01000011110011,
14'b00010011101110,
14'b00000010111110,
14'b00010010101010,
14'b00000110011101,
14'b00101000001100,
14'b00101111100011,
14'b00111110100000,
14'b00111100101011,
14'b00100110100011,
14'b00111010111011,
14'b00110100101110,
14'b00011010101110,
14'b00000000011011,
14'b00011010010110,
14'b00001101100111,
14'b00111100000111,
14'b00101001111100,
14'b00011101101001,
14'b00100000000100,
14'b00111111100001,
14'b00111110011101,
14'b00011111010111,
14'b00100010000001,
14'b00011001001000,
14'b00010000001110,
14'b00110000111101,
14'b00001010111011,
14'b00011111001100,
14'b00101111111000,
14'b01000000000101,
14'b00010101010101,
14'b00011011110001,
14'b01000001100100,
14'b00111101000011,
14'b00110110100000,
14'b00001110100011,
14'b00111000110110,
14'b00100001101100,
14'b00100100100100,
14'b00110011100001,
14'b00111110000101,
14'b00110011100101,
14'b00101000000100,
14'b00110111100000,
14'b00111110011011,
14'b00100011110010,
14'b00110010111110,
14'b00000010010111,
14'b00100000011001,
14'b00111100111010,
14'b00010011101100,
14'b00011111110000,
14'b00000010101100,
14'b00100010110000,
14'b00100101000110,
14'b00101001101111,
14'b00010101000010,
14'b00110111010001,
14'b00011010110001,
14'b00001110011000,
14'b00011000110000,
14'b00101100111010,
14'b00100101110000,
14'b00001111101011,
14'b00110110100011,
14'b00001011001001,
14'b00110111011000,
14'b00001110110000,
14'b00111110111110,
14'b00110010100101,
14'b00011001010011,
14'b01000000111110,
14'b00010010010101,
14'b00011110111000,
14'b00000111100100,
14'b00101001101011,
14'b00110111111011,
14'b01000101011011,
14'b00000111011101,
14'b01000010110111,
14'b00001100011010,
14'b00100100100000,
14'b00101000010010,
14'b00100111111011,
14'b00001001101111,
14'b00101001100101,
14'b00100010011100,
14'b00000001000001,
14'b00001010111000,
14'b00100111001101,
14'b00100001100010,
14'b00010100101000,
14'b01000011111001,
14'b01000000111000,
14'b00001110010011,
14'b00000101110000,
14'b00010110011010,
14'b01000010111001,
14'b00101001010100,
14'b00100011100010,
14'b00010101111000,
14'b00111100100000,
14'b00001010110011,
14'b00110001111000,
14'b00001010000100,
14'b01000110001011,
14'b00110101001101,
14'b01000111100000,
14'b00101000110011,
14'b00001010001110,
14'b00011010011110,
14'b00111000001000,
14'b00100000011010,
14'b00011001111001,
14'b00100110011010,
14'b01000101100000,
14'b00100101000001,
14'b00100000010101,
14'b00010100111100,
14'b00010101101010,
14'b00001111111011,
14'b00110010101001,
14'b01000000111011,
14'b00110111011001,
14'b00100010011110,
14'b00101100001001,
14'b00101111000011,
14'b00110001011000,
14'b00110000000001,
14'b01000100101000,
14'b00111011101011,
14'b00001111101010,
14'b00001100010111,
14'b00111111110101,
14'b01000101111101,
14'b00110010101010,
14'b00010010001001,
14'b00011101001110,
14'b01000010110101,
14'b00100001111010,
14'b00100101001111,
14'b00111011000000,
14'b00111001011111,
14'b00001100010100,
14'b00100111110000,
14'b00001001010001,
14'b00101010011010,
14'b01000001111001,
14'b01000011111010,
14'b00010101001001,
14'b00001011001110,
14'b00000000111111,
14'b00111000111000,
14'b00011011001000,
14'b00100011100101,
14'b00111010110010,
14'b00000010001011,
14'b00110100100000,
14'b00011111000111,
14'b00000110100001,
14'b00101100011110,
14'b00000111100011,
14'b00001101100011,
14'b00000111111001,
14'b01000110100001,
14'b00001111110111,
14'b00000010110111,
14'b00110001000110,
14'b00010101011110,
14'b00111011001001,
14'b00101000101101,
14'b00100111110001,
14'b00101101000100,
14'b00010111110010,
14'b00110101010011,
14'b00111000110101,
14'b00010000000001,
14'b00000101110001,
14'b00100001100001,
14'b00111100001010,
14'b00111110010000,
14'b00000100010001,
14'b00110011111001,
14'b01000101001111,
14'b01000100111100,
14'b00001010100001,
14'b01000001000111,
14'b00010010110011,
14'b00111111010000,
14'b01000100011000,
14'b00100101010001,
14'b00000101010111,
14'b00001001100001,
14'b00111010001110,
14'b00110111010100,
14'b00111100100100,
14'b00101100001011,
14'b00001101000000,
14'b00111110100110,
14'b01000000010100,
14'b00100001001111,
14'b00000111011110,
14'b00011100111110,
14'b00111100000000,
14'b00100010100011,
14'b00101111111101,
14'b00010001001111,
14'b01000010011111,
14'b00101010010101,
14'b00011001111010,
14'b01000001110111,
14'b00110100110010,
14'b00111111111010,
14'b00010110111111,
14'b01000000100010,
14'b00010100111000,
14'b00100000100011,
14'b00001100110101,
14'b00101011101111,
14'b00111010000000,
14'b00001011001000,
14'b00000110101011,
14'b00101110100110,
14'b00010000010010,
14'b00011010010010,
14'b00011101010110,
14'b00011101000100,
14'b01000110000100,
14'b00100001111100,
14'b00011100111010,
14'b00001001110111,
14'b00001001110100,
14'b00011001000010,
14'b00111111111011,
14'b00010110110101,
14'b00110101110101,
14'b00111000011000,
14'b00101111101101,
14'b00001110010010,
14'b00111010100110,
14'b00011100110000,
14'b01000101110000,
14'b00000010010100,
14'b00000110110011,
14'b00010111100000,
14'b00011101000010,
14'b00110011001010,
14'b01000111101100,
14'b01000100000111,
14'b00111101011111,
14'b00010100001000,
14'b00011101110100,
14'b00100000101011,
14'b00010000011010,
14'b00010010110101,
14'b00010001101010,
14'b00000000100111,
14'b00000000111000,
14'b00101110000010,
14'b01000100100011,
14'b00000110011000,
14'b00011010001111,
14'b00011011000010,
14'b00111011100010,
14'b00000110001011,
14'b00010000100010,
14'b00111111001111,
14'b00011110011110,
14'b00110001010010,
14'b00001011010001,
14'b00000001100010,
14'b00100110001111,
14'b00111111101001,
14'b00011110011000,
14'b00011000000000,
14'b00111001110001,
14'b00101011111001,
14'b00111000000111,
14'b00000010011110,
14'b00100010000011,
14'b00010010000010,
14'b00111110001000,
14'b00110001010111,
14'b00010001001010,
14'b00100110010111,
14'b00001100101001,
14'b00010000001000,
14'b00011110000010,
14'b00011001011000,
14'b00110100000001,
14'b00011010111101,
14'b01000000010000,
14'b00010110101001,
14'b00100010111100,
14'b01000011001101,
14'b00001111100110,
14'b00111000011010,
14'b00111110010111,
14'b00101001011111,
14'b00000011100110,
14'b00001010010110,
14'b00000011010010,
14'b00111100010011,
14'b00010010100110,
14'b00010101011011,
14'b00000000111101,
14'b00101000011110,
14'b00011000010110,
14'b00010001110100,
14'b00011110001001,
14'b00110110011100,
14'b00011100110100,
14'b00100110000010,
14'b00010110001001,
14'b00010001010010,
14'b00110111010011,
14'b00110000100101,
14'b00011110010011,
14'b00010000000110,
14'b00111001100110,
14'b00100011010001,
14'b00001000101010,
14'b01000101010100,
14'b00010110111000,
14'b00010000101111,
14'b00111111110001,
14'b00111100010010,
14'b00111101100111,
14'b00110011111011,
14'b00011000010000,
14'b00111011000001,
14'b00001110110111,
14'b00000000100011,
14'b00111100100110,
14'b00111111000111,
14'b00101001111110,
14'b00100000110000,
14'b00001100101100,
14'b00100011001010,
14'b00010001100100,
14'b00011110001101,
14'b00110110100001,
14'b00011101011001,
14'b00110000001010,
14'b01000010011100,
14'b00110111111101,
14'b00000111010111,
14'b00101000001110,
14'b01000001011010,
14'b00001111101111,
14'b00000111000100,
14'b00100110111011,
14'b00111100011101,
14'b00001111110001,
14'b00111010100101,
14'b00001101010111,
14'b00010111110110,
14'b00000110000010,
14'b00011000101001,
14'b00110010100110,
14'b00010100011110,
14'b00010110010110,
14'b00101111001101,
14'b00010101001101,
14'b00100100001110,
14'b01000100010000,
14'b00011010101101,
14'b00010100101100,
14'b00101011011001,
14'b00110001001011,
14'b00101001101110,
14'b00001010110100,
14'b01000101101111,
14'b00001101011111,
14'b00110101101100,
14'b01000011101101,
14'b00100000001101,
14'b01000000100110,
14'b00110011101010,
14'b00111100111110,
14'b00000000011101,
14'b00000101111100,
14'b00010101001100,
14'b00010100110000,
14'b00100110100110,
14'b00010100101111,
14'b00011101110000,
14'b00110100100101,
14'b00110011101111,
14'b00101100110001,
14'b00001111001011,
14'b00111010111111,
14'b00100101001010,
14'b00011000001010,
14'b00011111000110,
14'b00001110100110,
14'b00111100101101,
14'b00101101001001,
14'b00110100110101,
14'b00011101101000,
14'b00000011100011,
14'b00110110000111,
14'b00000110110111,
14'b00000111001011,
14'b00101011111100,
14'b01000011110110,
14'b00001010111100,
14'b00001110001110,
14'b00010100001110,
14'b00110010010100,
14'b00010110001011,
14'b00000101100111,
14'b00110111110011,
14'b00110110101000,
14'b00010111000011,
14'b00001000011000,
14'b00011001001100,
14'b00101100100111,
14'b00111111011011,
14'b00010010100000,
14'b00010101001111,
14'b00000101110010,
14'b00010010111110,
14'b00000101000100,
14'b00100001010000,
14'b00100000110101,
14'b00100101101011,
14'b00100000001001,
14'b00010100010011,
14'b00110001000000,
14'b00111111111111,
14'b00010010100011,
14'b00100000100001,
14'b01000110111100,
14'b00010010100001,
14'b00011001011100,
14'b00100110110100,
14'b00110100111100,
14'b00100010010010,
14'b00010000011111,
14'b00001101101010,
14'b00011101000001,
14'b00011110000001,
14'b00110001110111,
14'b00110100111010,
14'b00010010101111,
14'b01000100101011,
14'b00001001000100,
14'b00110101100110,
14'b00101000000101,
14'b00011011011010,
14'b00101001000010,
14'b00100001010011,
14'b01000100111101,
14'b00100110000101,
14'b00101010000111,
14'b00111111111000,
14'b00011001100001,
14'b00010011010100,
14'b00100001110010,
14'b00001001001100,
14'b00011101001010,
14'b00000000101001,
14'b00011111011111,
14'b00010010101000,
14'b00100100101001,
14'b01000100111110,
14'b00011011100110,
14'b00101010101011,
14'b00100010010100,
14'b00001010010101,
14'b00001110100111,
14'b00010101001010,
14'b00100010100001,
14'b00110001100000,
14'b00110101000100,
14'b01000110101100,
14'b00110011101011,
14'b00000011101100,
14'b00011000000111,
14'b01000111110111,
14'b00110101100100,
14'b00101010000100,
14'b00101111000000,
14'b00111011000110,
14'b00110100010100,
14'b00110111111111,
14'b00010101111110,
14'b01000010000110,
14'b00000110000110,
14'b00111000001110,
14'b00011100011110,
14'b00100111011000,
14'b01000111110010,
14'b00001011100101,
14'b00000001110111,
14'b00001111110011,
14'b00000100010100,
14'b00100000100010,
14'b00001110011100,
14'b00100010011101,
14'b00110100010111,
14'b00000000010100,
14'b00110110101010,
14'b00110010100010,
14'b00101000100011,
14'b00101011000100,
14'b01000111001110,
14'b00001010000110,
14'b00101000100001,
14'b00000011110100,
14'b00000100011000,
14'b00010011110010,
14'b00111110010110,
14'b01000010100010,
14'b00111000011011,
14'b00011000011011,
14'b00010100001010,
14'b01000101110010,
14'b00100010111110,
14'b00000101011011,
14'b00000010011000,
14'b00011011011001,
14'b00100100101110,
14'b00001100011100,
14'b00011010001001,
14'b00110010001111,
14'b00100011000011,
14'b00111010011100,
14'b00000111101110,
14'b01000000101011,
14'b00011001001011,
14'b00010011001111,
14'b01000100110001,
14'b00101001010001,
14'b00001111110110,
14'b00100101000011,
14'b00111001010000,
14'b00101011111101,
14'b00011011100011,
14'b00001011000000,
14'b00110111110001,
14'b00001111110010,
14'b00100110111001,
14'b00001001111011,
14'b00000110010101,
14'b00000101101101,
14'b00010101101101,
14'b00101001110010,
14'b00100110100101,
14'b01000011101010,
14'b00010110011000,
14'b00000111101010,
14'b00101000100100,
14'b00111011000010,
14'b00010010111100,
14'b00111011100111,
14'b00101000001101,
14'b00111010101011,
14'b00100010101111,
14'b00111001111000,
14'b00101110011101,
14'b00011111001111,
14'b00111111100110,
14'b00101110101101,
14'b00100111110010,
14'b00101000000000,
14'b00000111000011,
14'b00010111010000,
14'b01000110111011,
14'b01000100010011,
14'b00000010101110,
14'b00011001000000,
14'b00110000000100,
14'b00110011111010,
14'b00110010001110,
14'b01000001101000,
14'b00110000101001,
14'b01000000011111,
14'b00000100111001,
14'b00111101100011,
14'b00001101010100,
14'b00010000011110,
14'b01000111101011,
14'b00110100000010,
14'b00100010000010,
14'b00100000001010,
14'b00110101111111,
14'b00101100110111,
14'b00010001111100,
14'b00101110101010,
14'b00001000011111,
14'b00011000000011,
14'b00110000001110,
14'b00000111010011,
14'b00000010000000,
14'b00101011101010,
14'b00111000001001,
14'b00000011001110,
14'b00000110000100,
14'b00011001001001,
14'b00010011100001,
14'b00010011010110,
14'b01000111010011,
14'b00011110101010,
14'b00001010001101,
14'b00101011110000,
14'b01000011101100,
14'b00111010000010,
14'b01000001000001,
14'b00110011110010,
14'b01000110111110,
14'b00000011100101,
14'b00011000011111,
14'b00100111000111,
14'b01000011100001,
14'b00010011010101,
14'b00011000110101,
14'b00000000010111,
14'b00110010001000,
14'b00001101011001,
14'b00000000001010,
14'b00011000110110,
14'b00010000110000,
14'b00011000111011,
14'b00011010110000,
14'b00100100010101,
14'b00011100110011,
14'b00011010110011,
14'b00011011110000,
14'b01000100001000,
14'b00111101100001,
14'b00010110101101,
14'b00101001111101,
14'b00001101110101,
14'b00001010101001,
14'b00010100101110,
14'b00110010000001,
14'b00001001001110,
14'b01000010100110,
14'b00001000101101,
14'b00000001000010,
14'b00101010101110,
14'b00111010101100,
14'b00110011111110,
14'b00111100100101,
14'b00000011001000,
14'b00011011011110,
14'b00011110100110,
14'b00000100000110,
14'b00101000010011,
14'b00001110100010,
14'b00101110101001,
14'b00000110110101,
14'b00100110010000,
14'b00101001001010,
14'b00101111010110,
14'b00101011011010,
14'b01000110100011,
14'b00110100010010,
14'b00011111110011,
14'b00011100100011,
14'b01000110010010,
14'b00100000000001,
14'b01000101010001,
14'b00010110010001,
14'b01000111100111,
14'b00111011100001,
14'b00111110101001,
14'b00110111001110,
14'b00010110000010,
14'b00001010100111,
14'b00000100110101,
14'b00111101110001,
14'b00100111101101,
14'b00001010001010,
14'b00111001100001,
14'b00111001011011,
14'b00011000100110,
14'b01000001100010,
14'b00100110011100,
14'b00010011011011,
14'b00111110111100,
14'b00010110110110,
14'b00000000110010,
14'b00000001110000,
14'b00000110100010,
14'b00100111111001,
14'b00110101111001,
14'b01000001101001,
14'b00110110110100,
14'b00111001010111,
14'b00000110010110,
14'b00111111110100,
14'b00001101101000,
14'b00000000001100,
14'b00001001110001,
14'b00011100010000,
14'b00010101000001,
14'b00110010010011,
14'b01000111101000,
14'b00000000101101,
14'b00101010010010,
14'b00111110100010,
14'b00001001101010,
14'b00101111000001,
14'b00111011101100,
14'b00000100001000,
14'b01000011111101,
14'b00010100100110,
14'b00100001111101,
14'b00111101010100,
14'b00000011011101,
14'b00100100000100,
14'b00011010101000,
14'b00100111101010,
14'b00001000110001,
14'b00110110111110,
14'b01000000010101,
14'b00111110101110,
14'b00011100001011,
14'b00100010011000,
14'b00001010110001,
14'b00011000110100,
14'b01000001111010,
14'b00100101000000,
14'b00111111101011,
14'b00001101011000,
14'b00000101100101,
14'b00100000101010,
14'b00011000111100,
14'b00111010000100,
14'b00111010010111,
14'b00000011111111,
14'b00101011100110,
14'b00010100011010,
14'b00111100000011,
14'b00111110111001,
14'b00101000101110,
14'b00111111001000,
14'b00110100000111,
14'b00100000001011,
14'b01000000000111,
14'b00101000101100,
14'b00011101000111,
14'b00000000101010,
14'b00010111101111,
14'b00100100011101,
14'b00010010110111,
14'b00111001011010,
14'b00001000111100,
14'b01000110110111,
14'b00111000111010,
14'b00101111110001,
14'b00111000011101,
14'b00011001000011,
14'b00111001000010,
14'b00100100000001,
14'b00010111000101,
14'b00111000101101,
14'b00001000010101,
14'b00101111001000,
14'b00111011001100,
14'b00011010000000,
14'b00101110100101,
14'b00111110111010,
14'b00101011001000,
14'b00111001101100,
14'b01000011000110,
14'b00010101101111,
14'b01000010101100,
14'b00100111110100,
14'b00000001001010,
14'b00110011110011,
14'b00101111010010,
14'b00010110011100,
14'b00111001010001,
14'b00100000101000,
14'b00111110101000,
14'b00010000101110,
14'b00000100010110,
14'b00100100010100,
14'b00010001101100,
14'b00100101110011,
14'b00011001010010,
14'b00111010111001,
14'b00011010100110,
14'b00110001110101,
14'b00011011001010,
14'b00001111001110,
14'b00010010000110,
14'b00101001100110,
14'b00000011000101,
14'b00000001111100,
14'b00101011100001,
14'b00000011011010,
14'b00001111010001,
14'b00001101110011,
14'b00000001011100,
14'b00111111110000,
14'b00000110001001,
14'b00111110011000,
14'b00101001001101,
14'b00001101100001,
14'b00000011111100,
14'b00101010011101,
14'b00100110001101,
14'b00110000110000,
14'b00000010100100,
14'b00010000000000,
14'b00011111011101,
14'b00010010101101,
14'b00101110001010,
14'b00110101100101,
14'b00000000110111,
14'b00111010000101,
14'b00011101001111,
14'b01000110010111,
14'b00001001100011,
14'b00010111111110,
14'b00001111011000,
14'b00100110001000,
14'b00000001101111,
14'b00110011111100,
14'b00101011111111,
14'b00101100001100,
14'b01000001010110,
14'b00011101101111,
14'b01000001011100,
14'b00000101000010,
14'b00111011111000,
14'b00110111000101,
14'b00000111101101,
14'b00001000100011,
14'b00110011001011,
14'b00010100100101,
14'b00011111011010,
14'b00111001111010,
14'b00001111111111,
14'b00000001101100,
14'b00010001010110,
14'b00111010100100,
14'b00010011010011,
14'b00000111010101,
14'b00011010100101,
14'b01000110101110,
14'b00000110001100,
14'b00110000110111,
14'b00011010000101,
14'b00110101101110,
14'b00000100101010,
14'b00011100000110,
14'b00110011101000,
14'b01000010001000,
14'b00101111010111,
14'b00001000010011,
14'b00101100110010,
14'b00101001011100,
14'b01000100001100,
14'b00101000001001,
14'b00100100001000,
14'b00100010110101,
14'b01000111011111,
14'b00011000100101,
14'b00000110010000,
14'b00100010000100,
14'b00001101100100,
14'b01000110011000,
14'b00100000010110,
14'b00010010101011,
14'b00011011011101,
14'b00101100111101,
14'b00011100001110,
14'b00110110011001,
14'b00011101111000,
14'b00011100011010,
14'b00100101010101,
14'b00010010000001,
14'b00011011010011,
14'b00000011001111,
14'b01000100100101,
14'b00000111001000,
14'b00100110011001,
14'b01000110010101,
14'b00110001001001,
14'b00010110000011,
14'b00110010110101,
14'b00000100010111,
14'b00110001111011,
14'b00011101001011,
14'b00110011111000,
14'b00110010100000,
14'b00000011000010,
14'b00001100101101,
14'b00101111011110,
14'b00110100100011,
14'b00011110110010,
14'b00001101001100,
14'b00011000110111,
14'b00010100001101,
14'b00011011000011,
14'b00001001001111,
14'b00011111101100,
14'b01000101111100,
14'b00111101101101,
14'b00010111001000,
14'b00110101010010,
14'b00001001010111,
14'b01000100100110,
14'b00100010011001,
14'b00000110110110,
14'b00110111110111,
14'b00000110101100,
14'b00110110000100,
14'b00000100100001,
14'b00101101011011,
14'b00001100000100,
14'b00001011101000,
14'b01000110001111,
14'b00011011110011,
14'b01000110100111,
14'b00000100001011,
14'b00101011011110,
14'b00001010011010,
14'b00110000100001,
14'b00110100111101,
14'b00001011000111,
14'b00101010010000,
14'b00101001000101,
14'b00011111100000,
14'b00000111100001,
14'b00111010111000,
14'b00000000000100,
14'b00111001100000,
14'b00010001110001,
14'b00010011010010,
14'b01000101111011,
14'b00011111111011,
14'b00111100111101,
14'b00110111011101,
14'b00010011110011,
14'b00011010010111,
14'b00100111010110,
14'b00101101110110,
14'b00001101111100,
14'b00101000110001,
14'b00001101001011,
14'b00101001000111,
14'b00000000110101,
14'b00110000001001,
14'b00100110111110,
14'b00100000001111,
14'b00001100001101,
14'b00011100011001,
14'b00000100111111,
14'b00011111000001,
14'b00001010001111,
14'b00001011100111,
14'b00000010111111,
14'b00110101011000,
14'b00100001110000,
14'b00111111011101,
14'b00010111011001,
14'b00010110100110,
14'b00110010110011,
14'b01000110110110,
14'b00001110100100,
14'b00101011101011,
14'b00010110101100,
14'b00001101000110,
14'b00100111110110,
14'b00010011011001,
14'b00011101100011,
14'b00111110000100,
14'b00010110010100,
14'b00100010001000,
14'b00101000110101,
14'b00011000000101,
14'b00110111111010,
14'b00111100110010,
14'b00110000111110,
14'b00101011111000,
14'b00111011000101,
14'b00101101111111,
14'b01000001110011,
14'b00010011100100,
14'b00010001100011,
14'b00101010100111,
14'b00101111111111,
14'b00111011000111,
14'b00110001110100,
14'b01000000101111,
14'b00101001100010,
14'b00011001000110,
14'b00100001000101,
14'b00001101010010,
14'b00001001101101,
14'b00010101111101,
14'b00011100100100,
14'b00000110100000,
14'b01000000101000,
14'b01000110001100,
14'b01000000000001,
14'b00010001110011,
14'b00101011010010,
14'b00101110000000,
14'b00000110010001,
14'b00100001101010,
14'b00001000000011,
14'b00000111110000,
14'b01000011001110,
14'b00001100110111,
14'b00101011010000,
14'b00010100110100,
14'b00100100010111,
14'b00101110100000,
14'b01000101000001,
14'b01000001111000,
14'b00100100100011,
14'b00010011001110,
14'b00101110001111,
14'b00011010100000,
14'b00000111110110,
14'b00011100000001,
14'b00100110000011,
14'b01000001011011,
14'b00101011101000,
14'b00101111010011,
14'b01000011001010,
14'b00001110111101,
14'b00010000111001,
14'b00111000000001,
14'b01000010011101,
14'b00100001101001,
14'b00100100101111,
14'b00000100100110,
14'b00100110111010,
14'b00011111111101,
14'b00100111100110,
14'b00000110001110,
14'b00000010110010,
14'b00100011100001,
14'b00000101100100,
14'b00000100110110,
14'b00010101100001,
14'b00010111011000,
14'b00110010111100,
14'b00011100110101,
14'b00100110100001,
14'b00010101000100,
14'b00110110001011,
14'b01000111000110,
14'b00101011001100,
14'b00010111111010,
14'b00010011101111,
14'b01000000111010,
14'b00000101001100,
14'b00001011110011,
14'b00011001000100,
14'b00110100111111,
14'b00011010101011,
14'b00110111101111,
14'b01000010100111,
14'b01000111111001,
14'b01000010001110,
14'b00110010010001,
14'b00010011000000,
14'b00100000101001,
14'b00000011001011,
14'b00010110011111,
14'b00000010101111,
14'b00101010011001,
14'b00000010000101,
14'b00100011111011,
14'b00000001010110,
14'b00111100101110,
14'b00011101011010,
14'b00101010010111,
14'b00101010110001,
14'b00111000000011,
14'b00011111011001,
14'b00111010100000,
14'b00100100011011,
14'b00000100110010,
14'b00110110111001,
14'b00011001001010,
14'b00000001101010,
14'b00000101100011,
14'b00100101100101,
14'b00110010000000,
14'b00100010101001,
14'b00111110110011,
14'b00000000011001,
14'b00111011100100,
14'b00011101001001,
14'b01000011001011,
14'b00011010000111,
14'b00100001011100,
14'b00101000011000,
14'b00010100000010,
14'b00101100011101,
14'b01000101110001,
14'b00110011001100,
14'b00110101100111,
14'b00010001001011,
14'b00100101110100,
14'b00110001111001,
14'b00101000001111,
14'b00000111110001,
14'b00000111111000,
14'b00111001001000,
14'b01000111010111,
14'b00011110110111,
14'b00010010111011,
14'b00000110011100,
14'b00011110100100,
14'b00110101101011,
14'b00111111001010,
14'b00001101000111,
14'b00100011000001,
14'b00101000101111,
14'b00011010111100,
14'b00000000000001,
14'b00000101010101,
14'b01000111010101,
14'b00010101010000,
14'b00101101100100,
14'b00100111011101,
14'b00010001000000,
14'b00101010011011,
14'b00010100000111,
14'b00000101000110,
14'b00000001100011,
14'b00111011100000,
14'b00011011010111,
14'b00000001010010,
14'b00101000111000,
14'b00000101011010,
14'b00011001100111,
14'b01000000100000,
14'b00101111000101,
14'b00100010101101,
14'b00111110001111,
14'b00001000010001,
14'b00100001101000,
14'b00010010010011,
14'b00001011111011,
14'b00100100000110,
14'b00011110000110,
14'b00001101010011,
14'b00100010001111,
14'b00010100000001,
14'b00000100110011,
14'b00111100001001,
14'b00000000100110,
14'b00101010110000,
14'b00000110111110,
14'b00000000010010,
14'b00111100110111,
14'b00100100001010,
14'b00010001111000,
14'b00100000010011,
14'b00001100000000,
14'b00010010010111,
14'b00010110100101,
14'b00011011101011,
14'b00010111011110,
14'b00101011001111,
14'b00011000100100,
14'b00001101001110,
14'b01000011101011,
14'b00101011000101,
14'b00001010110111,
14'b00110011110101,
14'b01000011110001,
14'b00111100000101,
14'b01000000111100,
14'b00001010100011,
14'b00110111111000,
14'b00001000110101,
14'b00100000011011,
14'b00100000000101,
14'b00001010100110,
14'b00111010010110,
14'b00101001111111,
14'b00010100101010,
14'b00001001111000,
14'b00010111000100,
14'b00011100001000,
14'b01000000001100,
14'b00001111101100,
14'b00011111110010,
14'b00011111010100,
14'b00000111011100,
14'b00011010011001,
14'b01000110010001,
14'b00101100100110,
14'b00000011110001,
14'b00011011100101,
14'b01000000110111,
14'b00001111000000,
14'b01000101001101,
14'b00010110101010,
14'b00000100100010,
14'b01000101111010,
14'b00110001010100,
14'b00111101010000,
14'b00001011010011,
14'b00010101010100,
14'b00011100010001,
14'b00011100011111,
14'b00010111101110,
14'b00101101000001,
14'b01000111111101,
14'b00000101000000,
14'b00100010111101,
14'b00110100101100,
14'b00011001111011,
14'b00011110001000,
14'b01000011000100,
14'b00100110001001,
14'b00100100101100,
14'b00010000110110,
14'b00101110001001,
14'b00000001000000,
14'b00000101101010,
14'b01000110000011,
14'b00000101010011,
14'b00110010011100,
14'b00001100101000,
14'b00000101011000,
14'b00011000000001,
14'b00001110001000,
14'b00111111010010,
14'b00010101110000,
14'b01000101001001,
14'b00101111111011,
14'b00101110110101,
14'b00111110110001,
14'b00111101000111,
14'b00111111111100,
14'b00001011011011,
14'b00000100110000,
14'b00100001000011,
14'b00101011101110,
14'b00001011001011,
14'b00000011100001,
14'b00100111101001,
14'b00110011010110,
14'b00010111101011,
14'b00100000110110,
14'b00001101110111,
14'b00100101011110,
14'b00010001111011,
14'b00101011011100,
14'b00101100100100,
14'b00101001100000,
14'b00101100001111,
14'b00001111100101,
14'b00100111011011,
14'b01000110001001,
14'b00010010011000,
14'b00110001100110,
14'b00101001101000,
14'b00110110111111,
14'b00011011100000,
14'b00100110000000,
14'b00111001000101,
14'b00110001101111,
14'b00100001010010,
14'b00000011010000,
14'b00101001001001,
14'b00111000000010,
14'b00110000100100,
14'b00001100110100,
14'b01000100011011,
14'b01000101000100,
14'b00001110010001,
14'b01000011100100,
14'b00001011111000,
14'b00111010011001,
14'b00001011100000,
14'b00010101100101,
14'b00000000101111,
14'b00101101000111,
14'b01000110001000,
14'b00010010001100,
14'b00001110001100,
14'b00111100011111,
14'b00011011011111,
14'b00010000000111,
14'b01000110100000,
14'b00100010001110,
14'b00011100011000,
14'b00110101000011,
14'b00101011100000,
14'b00010000101101,
14'b00101111011001,
14'b00000000010000,
14'b00100000111110,
14'b01000101111000,
14'b01000110101010,
14'b00110000001111,
14'b00111001101000,
14'b00111001100011,
14'b01000100111001,
14'b01000001100000,
14'b00101000110000,
14'b00010000001111,
14'b00101011000000,
14'b00111100000110,
14'b00011000100000,
14'b00111101110100,
14'b00011101100110,
14'b00000111011111,
14'b00111111001110,
14'b01000011011100,
14'b00011000101111,
14'b00010001100111,
14'b00110000111100,
14'b00101111111110,
14'b00011110010100,
14'b00110111100110,
14'b00000001001011,
14'b00000011100111,
14'b00100000000110,
14'b00101111110111,
14'b00101000111111,
14'b00110010011110,
14'b00111010110000,
14'b00110110101011,
14'b00011001110000,
14'b00110001000100,
14'b00110000010101,
14'b00010001001101,
14'b00011110101011,
14'b00100000011111,
14'b00111011101010,
14'b00001110101110,
14'b01000001101010,
14'b00001001000001,
14'b00001100110010,
14'b00111111011010,
14'b00101110100100,
14'b00110000101110,
14'b00001011101111,
14'b00011101110010,
14'b00011110100010,
14'b00011011101110,
14'b00000101110110,
14'b00010110110100,
14'b01000011001100,
14'b00110111101010,
14'b00101110110001,
14'b01000101011001,
14'b00111001110101,
14'b00101001101010,
14'b00110011100111,
14'b00100001110110,
14'b00111110111011,
14'b00100101101010,
14'b00100011111101,
14'b00000110110000,
14'b00011100100111,
14'b00011110111010,
14'b00010011111010,
14'b00110010100100,
14'b01000111110101,
14'b00010000010110,
14'b00010000001010,
14'b00100011100100,
14'b00100100101010,
14'b00101110011000,
14'b00110001011101,
14'b00111000111101,
14'b00000100101001,
14'b01000010111010,
14'b00111110001110,
14'b00111101111010,
14'b00001100001010,
14'b00101101000000,
14'b00010001000110,
14'b00010100100111,
14'b00110101111011,
14'b00110000110001,
14'b00100011011111,
14'b00101101011100,
14'b00100110110011,
14'b00100011001100,
14'b00000011110010,
14'b01000000011100,
14'b01000010010100,
14'b00011010010000,
14'b00101110110110,
14'b00011000100010,
14'b00011101100000,
14'b00010110010111,
14'b00011010001011,
14'b00011001011101,
14'b00001011110000,
14'b00010001101111,
14'b00011110011001,
14'b00110111001111,
14'b00100111111110,
14'b01000010100100,
14'b01000010110001,
14'b00000111111100,
14'b00011101000011,
14'b00011100001100,
14'b00001001010101,
14'b00101101111110,
14'b00010010110001,
14'b00010111010100,
14'b00010001000100,
14'b00010000001100,
14'b00000011010011,
14'b00011100001010,
14'b00001100111000,
14'b00000101101110,
14'b01000110101011,
14'b00101010000110,
14'b00000101110111,
14'b00101010111100,
14'b00101011010110,
14'b01000001010000,
14'b00000110110100,
14'b00101001011101,
14'b00000011010001,
14'b00011101110001,
14'b00001011011110,
14'b00100101011001,
14'b00111010001111,
14'b01000011000000,
14'b00101010010001,
14'b00101010110101,
14'b00010100110011,
14'b00110110010000,
14'b00101111001100,
14'b00001011111101,
14'b00101110000101,
14'b00000110011110,
14'b00111000010001,
14'b00011010100010,
14'b00001110101010,
14'b00010001110111,
14'b00001111001101,
14'b00000110111001,
14'b01000011101000,
14'b00010100000000,
14'b00000101000111,
14'b00111001010011,
14'b00001101101001,
14'b00011010111000,
14'b00110011010000,
14'b00111001000110,
14'b00100011101001,
14'b00111110000010,
14'b00100111001100,
14'b00010100010001,
14'b00011111101011,
14'b00111110000110,
14'b00100100110110,
14'b00111100010001,
14'b00110010000010,
14'b00010001010100,
14'b00100110101100,
14'b00110100000100,
14'b00001110001101,
14'b00000111011000,
14'b00110101000101,
14'b00010001010001,
14'b00010000111110,
14'b00111110110010,
14'b00010110100010,
14'b00011001110111,
14'b00100101010000,
14'b00101100100001,
14'b00101011001001,
14'b00010001111111,
14'b00111101000110,
14'b00000100101111,
14'b00011100101101,
14'b01000010011011,
14'b00001100001001,
14'b00110101100000,
14'b00010000010100,
14'b00000011111110,
14'b00001100000001,
14'b00110100101000,
14'b00011111010011,
14'b00111101101100,
14'b00100101100110,
14'b00001000110111,
14'b00101101111011,
14'b00000001100001,
14'b01000111011010,
14'b00011001110011,
14'b00100000000011,
14'b00010011111001,
14'b00110110111011,
14'b00010010100010,
14'b00101100011100,
14'b00111101001010,
14'b00011110000000,
14'b00101001010111,
14'b00111000111110,
14'b00011101101101,
14'b00111010111010,
14'b00111111110010,
14'b00011001100000,
14'b00001010101000,
14'b00010111110100,
14'b00111000010010,
14'b00010101011101,
14'b00011100100000,
14'b01000111100110,
14'b00100011010111,
14'b00000001110101,
14'b00111111011000,
14'b00101101100111,
14'b00110110000110,
14'b00001011100100,
14'b00010101001011,
14'b00010010011100,
14'b00001010011100,
14'b00101011111010,
14'b00001010001100,
14'b00010000000100,
14'b01000111000100,
14'b01000100100111,
14'b00010001011000,
14'b00101001011110,
14'b00110000101111,
14'b00011011000110,
14'b00110100001111,
14'b00001011101100,
14'b01000001111100,
14'b00100010001011,
14'b00001111111101,
14'b00110001000111,
14'b00111111111101,
14'b00110110000001,
14'b00101101110101,
14'b00111010001011,
14'b00010100001001,
14'b01000011000010,
14'b00111111000000,
14'b00101001001100,
14'b00011101000110,
14'b00001111000011,
14'b00110111110000,
14'b00001011011000,
14'b00101110000011,
14'b00000000001101,
14'b00001010011001,
14'b00000111110010,
14'b00101101010010,
14'b00000001001000,
14'b00011000111001,
14'b00000100110001,
14'b00000001111011,
14'b00110110001110,
14'b00011001011110,
14'b00011010000110,
14'b00101010010100,
14'b00111010010011,
14'b00000001111110,
14'b00001100111101,
14'b00110111101101,
14'b00101111110010,
14'b01000111001101,
14'b00001001001000,
14'b00000000100101,
14'b00001011001111,
14'b01000001000011,
14'b00011111100011,
14'b00111001111110,
14'b01000000100101,
14'b00001011101110,
14'b00110101110100,
14'b00011111000101,
14'b00010001010111,
14'b00001010111111,
14'b00011010101001,
14'b00011011000000,
14'b00010011101011,
14'b00001110100001,
14'b00110110111010,
14'b00010000101001,
14'b01000011111110,
14'b00111100010111,
14'b00001111101101,
14'b01000001001100,
14'b00001100001000,
14'b00010000010001,
14'b00010100100011,
14'b00011111011000,
14'b00001110101101,
14'b00110000110101,
14'b01000000011010,
14'b00001100010001,
14'b00010000010011,
14'b00100110011000,
14'b01000011100010,
14'b00001101100110,
14'b00111000111011,
14'b00110101110000,
14'b00111011111010,
14'b00001000001110,
14'b00001100000110,
14'b00100110000100,
14'b00000001011111,
14'b00000101110100,
14'b01000111011101,
14'b00100000101111,
14'b00111010010010,
14'b00010111100110,
14'b00011010010100,
14'b00111001010101,
14'b00111101011100,
14'b00001110000000,
14'b01000000000000,
14'b01000110001101,
14'b00101010000000,
14'b00010010001110,
14'b00001110000101,
14'b00001000110000,
14'b00111011101110,
14'b00110101001100,
14'b01000001010101,
14'b00011011100001,
14'b00100111100000,
14'b00110001111100,
14'b00110101011111,
14'b00001110100101,
14'b00101100100010,
14'b00111110100011,
14'b00110100001100,
14'b00000110100110,
14'b00111101010101,
14'b00011010001000,
14'b00110010001101,
14'b00111100111100,
14'b00101111100110,
14'b00100001110100,
14'b00001110010110,
14'b00101100101001,
14'b00001001101100,
14'b00011110010101,
14'b00011001001110,
14'b00000000111110,
14'b00011101110110,
14'b00110111000100,
14'b00000100011011,
14'b00111111100000,
14'b00110100111011,
14'b00111001101111,
14'b01000011011111,
14'b00100001100011,
14'b00001001111100,
14'b00101111011111,
14'b00011101101110,
14'b00100110010101,
14'b00011001010001,
14'b00010110110111,
14'b01000010010101,
14'b01000000000110,
14'b00000100000111,
14'b00100101000101,
14'b00010001011110,
14'b00010101000101,
14'b00111000000000,
14'b00010000011100,
14'b00000000100000,
14'b00001010000000,
14'b00011100100010,
14'b00000110010010,
14'b00100111110011,
14'b00100111100001,
14'b00110111100111,
14'b00000100101011,
14'b00011100101100,
14'b00110100101010,
14'b00011011010001,
14'b00110110010100,
14'b00111100001111,
14'b00001000110110,
14'b00110011110110,
14'b00000100000101,
14'b00000000001111,
14'b00110000100000,
14'b00110010001100,
14'b01000010000000,
14'b01000000011011,
14'b00111111100010,
14'b00110000001101,
14'b00100111100101,
14'b00001000100010,
14'b00101011010100,
14'b00001000000000,
14'b00001111011100,
14'b01000011101001,
14'b00000011011111,
14'b00111111111110,
14'b00101001000110,
14'b01000000100011,
14'b00001001110110,
14'b01000011010001,
14'b00110110011010,
14'b00101011111011,
14'b00011100010100,
14'b00000001010101,
14'b00110011000111,
14'b00010000011101,
14'b00001110011111,
14'b00101010101111,
14'b00011101100111,
14'b00100000000010,
14'b00111000010011,
14'b00101110010000,
14'b00100011110100,
14'b00001001110011,
14'b00000110011111,
14'b00100010010011,
14'b00001011010010,
14'b01000010101111,
14'b00011111100111,
14'b00101111110000,
14'b00110100110110,
14'b00101101100000,
14'b00110000101011,
14'b00001100111011,
14'b00010010000011,
14'b00010001101000,
14'b00001110111001,
14'b00100101010111,
14'b00100010110010,
14'b00010100011111,
14'b00001001001101,
14'b00010000101100,
14'b00011000000010,
14'b01000000000100,
14'b00101101101011,
14'b00110001111111,
14'b00101110110000,
14'b00111001110100,
14'b00010010011101,
14'b00011000001000,
14'b00110000011001,
14'b00001100010000,
14'b00010011011010,
14'b00000000111100,
14'b01000111010010,
14'b00001010111010,
14'b00011110000111,
14'b00101010101101,
14'b01000101100100,
14'b01000000111101,
14'b00000100110111,
14'b00000000111011,
14'b00000001000111,
14'b00000010001001,
14'b00011110111100,
14'b00110011001110,
14'b00000000010110,
14'b00001111011001,
14'b01000111110110,
14'b00011011101101,
14'b00010101100110,
14'b00110110111101,
14'b00001000001100,
14'b00101101101110,
14'b00001000101111,
14'b00000011100010,
14'b00001001110000,
14'b00000010010001,
14'b00000110101111,
14'b00111100111011,
14'b00111011001111,
14'b00110001000010,
14'b00011101111101,
14'b00010001111010,
14'b00100001111111,
14'b00101011101001,
14'b00100011101111,
14'b00000110111011,
14'b00001001010110,
14'b00000101111000,
14'b00011101001000,
14'b00110100100100,
14'b00010010111001,
14'b00110001001000,
14'b00000010100011,
14'b01000101011101,
14'b00001100011011,
14'b00010000110100,
14'b00100010100110,
14'b00110101000010,
14'b00000010111001,
14'b00011000011010,
14'b00011011111111,
14'b00010010001101,
14'b00001011010111,
14'b00010001001000,
14'b00011000010001,
14'b00100111001010,
14'b00010111110101,
14'b00000011110000,
14'b00111101100100,
14'b00111101101110,
14'b00110011011001,
14'b01000000011001,
14'b00100011000111,
14'b00110010000100,
14'b00110101001111,
14'b00001000000100,
14'b00001100010011,
14'b00100010001001,
14'b00010110111010,
14'b00000011110111,
14'b00110100101101,
14'b00001000110010,
14'b00010000110001,
14'b00000001010111,
14'b00101101110011,
14'b00101110111100,
14'b00011101101011,
14'b00111101100000,
14'b00101101011101,
14'b00101111011101,
14'b00000000111001,
14'b00111101101010,
14'b00000000000010,
14'b00100101010010,
14'b00011111000011,
14'b00100111100010,
14'b00010000110101,
14'b00001000100001,
14'b00101110100111,
14'b00110011100000,
14'b00110000010010,
14'b00100100000000,
14'b00101010100101,
14'b00110011111111,
14'b00010110111011,
14'b01000001110110,
14'b00001011110010,
14'b00100100101000,
14'b00001011101010,
14'b00011111001000,
14'b00101011110101,
14'b00111101010010,
14'b01000011000101,
14'b00010100111011,
14'b00001001100000,
14'b00101011011000,
14'b00001101000011,
14'b00000100010011,
14'b00111000011110,
14'b00001001101011,
14'b00110110101110,
14'b00011111011011,
14'b00100011101000,
14'b00111110000011,
14'b00011110010000,
14'b00111110000001,
14'b00011110001011,
14'b00000110000101,
14'b00110000000110,
14'b01000001110010,
14'b00001011100010,
14'b01000100010001,
14'b00110111100010,
14'b00110001010001,
14'b00001010101111,
14'b00011011001111,
14'b00111101000000,
14'b00010001101110,
14'b01000000010001,
14'b00001001110010,
14'b00001100100111,
14'b00011011101100,
14'b00011000101101,
14'b00111011011100,
14'b00010011110110,
14'b00111000010110,
14'b01000001010010,
14'b00010000111101,
14'b00100100111101,
14'b00000110001000,
14'b00011010011000,
14'b01000100101101,
14'b00101011001101,
14'b00100010110001,
14'b00010001011111,
14'b00110001100100,
14'b00111010110001,
14'b01000101010101,
14'b00011110010001,
14'b00111011110110,
14'b00011111010110,
14'b00100101000100,
14'b00001000100000,
14'b00101001110100,
14'b00100001011010,
14'b00100101010011,
14'b00000001001001,
14'b00100111000010,
14'b01000011110101,
14'b00100111101011,
14'b00011101001101,
14'b00000001100110,
14'b00000101100010,
14'b00010011110111,
14'b00000001011011,
14'b00111001001110,
14'b00000111111010,
14'b00000010010101,
14'b00001100011111,
14'b00000010010011,
14'b00100001000111,
14'b00110110110011,
14'b01000000010110,
14'b00010011000100,
14'b00111111100111,
14'b00100011110101,
14'b00111101001100,
14'b00100111011010,
14'b01000011000011,
14'b00001001100101,
14'b00010111101010,
14'b00000110010100,
14'b00111000101001,
14'b00000001111010,
14'b00101011010001,
14'b00101101001101,
14'b01000110101101,
14'b00000101010100,
14'b00011110001100,
14'b00001111000101,
14'b01000010110011,
14'b00111001000001,
14'b00001100000101,
14'b00001011110110,
14'b00011001000101,
14'b00000111000010,
14'b00101100000110,
14'b00010110000101,
14'b00101101100010,
14'b00101100110110,
14'b00010010000111,
14'b00101001101001,
14'b00001111000001,
14'b00000100010101,
14'b00110100110000,
14'b00110101010110,
14'b00000011111101,
14'b00111011110100,
14'b00100000010000,
14'b01000001111110,
14'b00100010000110,
14'b00011011011011,
14'b00011101111011,
14'b00111001100101,
14'b00111001000100,
14'b00001111110101,
14'b00000110011001,
14'b00100111110101,
14'b01000110010000,
14'b00110011100010,
14'b00001001010011,
14'b00010111110111,
14'b00010001001001,
14'b00010000111011,
14'b00011000100001,
14'b00111011011001,
14'b00100011011001,
14'b00101101101001,
14'b00010011101001,
14'b00001001101000,
14'b00001101101101,
14'b00100101011101,
14'b00000101010000,
14'b01000110000001,
14'b00000010001111,
14'b00110110110000,
14'b00000110101010,
14'b01000101110111,
14'b00001011110100,
14'b00011100111001,
14'b01000101111111,
14'b01000110100110,
14'b00011110010110,
14'b00000010111101,
14'b00100010100111,
14'b00001110111011,
14'b00111001111101,
14'b00010011010000,
14'b00110101010000,
14'b00010110010000,
14'b00101111010001,
14'b00110001100111,
14'b00111111000010,
14'b01000110011111,
14'b00000111000101,
14'b00000101000101,
14'b00100100000010,
14'b00001010100101,
14'b00000001011110,
14'b00100010001100,
14'b00111000100001,
14'b00000110010011,
14'b00010001100101,
14'b00101001000000,
14'b00110010011000,
14'b00110010011111,
14'b00001111111110,
14'b00000101010010,
14'b00000000111010,
14'b00110110011111,
14'b00011111101111,
14'b00001110101111,
14'b00110010101110,
14'b00110100111000,
14'b00001000011011,
14'b00111001100100,
14'b01000100110011,
14'b00101100111001,
14'b00001010000001,
14'b00100001110111,
14'b00001000001011,
14'b00000010110110,
14'b00101101100101,
14'b00011100101001,
14'b00001010010001,
14'b00011000100011,
14'b00011101010011,
14'b00110111001101,
14'b00101111101011,
14'b00111001010010,
14'b00100011111100,
14'b00110010111011,
14'b01000010101010,
14'b00010001100010,
14'b01000101111001,
14'b00011100010111,
14'b01000110110101,
14'b00110110011011,
14'b00110011011011,
14'b00110111000011,
14'b00101111110011,
14'b00010111010001,
14'b00000101111011,
14'b00010101010010,
14'b00101101001010,
14'b00100100110010,
14'b00001100111001,
14'b00111100110100,
14'b01000001000101,
14'b00110110100110,
14'b01000111010100,
14'b00110100001010,
14'b00111010011010,
14'b00100011110011,
14'b01000110111111,
14'b01000101000000,
14'b00101101011010,
14'b01000100011010,
14'b00100110001110,
14'b01000000100111,
14'b00101000100000,
14'b00101011010101,
14'b01000110110000,
14'b00110001101001,
14'b00110111110101,
14'b00110110110101,
14'b00110001110000,
14'b00001010000111,
14'b00010000100001,
14'b01000000101110,
14'b00111011110000,
14'b00111100101010,
14'b00000100100100,
14'b00001000011101,
14'b00001101001010,
14'b01000011101110,
14'b00001000001101,
14'b00100011000100,
14'b00111011100011,
14'b00111100000010,
14'b00101010110111,
14'b00111000000100,
14'b00101101110010,
14'b01000101101000,
14'b00011011010110,
14'b00010110110011,
14'b00001111110100,
14'b00111110110000,
14'b00100001001010,
14'b01000110000111,
14'b01000010100101,
14'b00010001000101,
14'b00101110111011,
14'b00110110011101,
14'b00101000011010,
14'b00101101011110,
14'b00100011100011,
14'b00001101010001,
14'b00100000010001,
14'b00001010011110,
14'b00110110010011,
14'b00010000111100,
14'b00110111010110,
14'b00110010001010,
14'b00101100110011,
14'b00010101011001,
14'b00010101110100,
14'b00101110011111,
14'b00111011100110,
14'b01000101101001,
14'b00000101001010,
14'b00011000111010,
14'b00100001111110,
14'b00011101101010,
14'b00010100101011,
14'b00001011010110,
14'b00010100100001,
14'b00011111001001,
14'b00101001001011,
14'b01000001101100,
14'b00101000011001,
14'b00100011011110,
14'b00111100101001,
14'b00111011111111,
14'b00011100010110,
14'b00101100100101,
14'b00011011001100,
14'b00110000000101,
14'b01000101000101,
14'b00001001111110,
14'b00100010111111,
14'b00110011101100,
14'b00001111100000,
14'b01000001011101,
14'b00000010110011,
14'b00101010101000,
14'b00100100111001,
14'b00011011001110,
14'b00011011001011,
14'b00010011100011,
14'b00100100001011,
14'b01000001000000,
14'b00010111100010,
14'b01000110011100,
14'b00110001001101,
14'b00110011111101,
14'b00111111101110,
14'b00110011000000,
14'b00101110100010,
14'b00111111000110,
14'b00111011111101,
14'b00111010111100,
14'b00001101111110,
14'b00000100001001,
14'b00000000011010,
14'b00010011011100,
14'b00110010111111,
14'b00100111001000,
14'b00100000111000,
14'b00011110100011,
14'b00110010101101,
14'b00111001101110,
14'b01000111010001,
14'b00101101100011,
14'b00001011011010,
14'b00110000010110,
14'b00100010110011,
14'b00011011110111,
14'b01000111000010,
14'b00000111010000,
14'b00010010110010,
14'b00011101100001,
14'b00000111000111,
14'b00110101110111,
14'b00000001100111,
14'b00111010011111,
14'b00001100100101,
14'b00101111011100,
14'b01000100000011,
14'b00110000111111,
14'b00011010110010,
14'b01000100010010,
14'b00101100000000,
14'b00000111010100,
14'b00000001101110,
14'b00100001100110,
14'b00110010101100,
14'b00010010110110,
14'b00110111101011,
14'b00000100011100,
14'b00100101101110,
14'b00101111001001,
14'b00101111101110,
14'b00010100001100,
14'b00100010111010,
14'b00101010100110,
14'b00000100101100,
14'b01000001000010,
14'b00001001011110,
14'b00010011001100,
14'b00110001001110,
14'b00100000100101,
14'b00110010111000,
14'b00111001101011,
14'b00010101101011,
14'b00101100001010,
14'b00010010010110,
14'b00101001110111,
14'b00001110111100,
14'b00011111110111,
14'b00111011111011,
14'b00100000111111,
14'b00110011100011,
14'b00011010100011,
14'b00001000001111,
14'b00101001010010,
14'b00110100010011,
14'b00001001000000,
14'b00001010100000,
14'b00000011100000,
14'b00011110101001,
14'b01000001001011,
14'b00101111110110,
14'b00100100111110,
14'b00001100111111,
14'b00111000100010,
14'b01000101110110,
14'b00111011001010,
14'b00101110110010,
14'b00100110110000,
14'b00110110110001,
14'b00101101010110,
14'b00000011010110,
14'b00011100101111,
14'b00110010010111,
14'b00010001100110,
14'b00000010011100,
14'b00100110011110,
14'b00011000000110,
14'b00110011000100,
14'b00011111010000,
14'b00011011001101,
14'b00101010111110,
14'b00110011000001,
14'b00001110001011,
14'b00100100011100,
14'b00011111010010,
14'b00011101011011,
14'b00110110100010,
14'b00100100011001,
14'b00111011011010,
14'b00110000001000,
14'b00001001000011,
14'b00001101010110,
14'b00011010111011,
14'b01000000001110,
14'b00101011000001,
14'b00010000101011,
14'b00110001111010,
14'b00111000001111,
14'b00000111010001,
14'b00101010010011,
14'b00011100011101,
14'b00110001100001,
14'b00010100111001,
14'b01000101001000,
14'b00111000110000,
14'b00101101110111,
14'b00111000100000,
14'b00000111000000,
14'b00111010000001,
14'b01000100101111,
14'b00111001111100,
14'b00100111101110,
14'b00110111011011,
14'b00101101001011,
14'b01000010101110,
14'b00001010011101,
14'b00100110101011,
14'b00111110111000,
14'b00111010001000,
14'b00101011001010,
14'b00010001010000,
14'b00110000101101,
14'b00111110101100,
14'b00010101011010,
14'b01000010000100,
14'b00011100001101,
14'b00101000011100,
14'b01000001100011,
14'b00111000001010,
14'b00101000100111,
14'b00110110010001,
14'b00001000101011,
14'b01000000001010,
14'b00111100010100,
14'b00011000001111,
14'b00110000010001,
14'b00001110110101,
14'b00010101000011,
14'b00101011001011,
14'b01000101100101,
14'b01000000101001,
14'b00001010110010,
14'b00001101111010,
14'b00001100010101,
14'b00010110100011,
14'b00000011101010,
14'b00110100011011,
14'b00100010010001,
14'b01000111101111,
14'b00101000101000,
14'b00101011100101,
14'b00111011110001,
14'b00011111100001,
14'b00111010111110,
14'b01000100011100,
14'b01000001010100,
14'b01000010000101,
14'b00100011110111,
14'b00101000111001,
14'b01000000101100,
14'b00011101111100,
14'b00011010010101,
14'b01000111001010,
14'b00110101010100,
14'b00101010111010,
14'b00100010100100,
14'b00011011100100,
14'b00101010001000,
14'b00001111011110,
14'b00000101101001,
14'b00001100001111,
14'b00101111000100,
14'b01000010001011,
14'b00111011101001,
14'b00010111010101,
14'b00111110111111,
14'b00100000001100,
14'b00110000101000,
14'b00100001011011,
14'b00011110000100,
14'b01000110011010,
14'b01000101101100,
14'b00001001100111,
14'b00110000001011,
14'b00000111001010,
14'b00111001110111,
14'b00111110001010,
14'b00001110011110,
14'b00000101000001,
14'b00011111001010,
14'b00001000111110,
14'b01000100001101,
14'b00110010101000,
14'b00110000001100,
14'b00001011000011,
14'b00010111010010,
14'b00110011010010,
14'b00110001001100,
14'b00101001111010,
14'b00011001010111,
14'b00011101001100,
14'b00011100110111,
14'b01000110111000,
14'b00101110010100,
14'b00100001010110,
14'b00101001100001,
14'b00100100100010,
14'b00001110011101,
14'b01000001100111,
14'b00110110100101,
14'b00000010100001,
14'b00111111101000,
14'b00100011000101,
14'b00000100000010,
14'b00110110011000,
14'b00101100101000,
14'b00100101001000,
14'b00110111110100,
14'b00001101100101,
14'b01000001000110,
14'b00010011000011,
14'b00000011000011,
14'b00110101011011,
14'b00100100000101,
14'b01000110000110,
14'b00110111000110,
14'b01000101010011,
14'b00000010101010,
14'b00011010001010,
14'b00100111100111,
14'b00100100001100,
14'b00101010110110,
14'b00110001011110,
14'b01000101101011,
14'b00111011110101,
14'b01000010111110,
14'b00110111000111,
14'b00000010100110,
14'b01000110101111,
14'b00110110101101,
14'b00000111100101,
14'b00101101111100,
14'b00100000100000,
14'b00010001101011,
14'b00111011110010,
14'b00011100111100,
14'b01000111101001,
14'b00000010110001,
14'b00111110101111,
14'b00000010000110,
14'b00010011111000,
14'b01000111010000,
14'b00001110110011,
14'b01000100001111,
14'b00101101010001,
14'b00100011001001,
14'b00100001001110,
14'b00000111110100,
14'b01000001100101,
14'b01000000110001,
14'b00000001011010,
14'b00000111011011,
14'b00111101110011,
14'b00011010011100,
14'b00101000101010,
14'b00000010111010,
14'b00110101011101,
14'b00000010010010,
14'b00100011001110,
14'b00100100101101,
14'b00000001011101,
14'b00000111011010,
14'b01000111001100,
14'b00110100111110,
14'b00010110110010,
14'b00111111010100,
14'b00001000010100,
14'b00000111101011,
14'b00101000010110,
14'b00100100100110,
14'b00011001111111,
14'b00001111101110,
14'b00110111111001,
14'b00001000111011,
14'b00001110011001,
14'b00100100010011,
14'b00000000100010,
14'b00110110101111,
14'b00001100110110,
14'b00101101011001,
14'b00100111111000,
14'b00010000000101,
14'b00011110110101,
14'b00010011011110,
14'b01000011010110,
14'b00101000110010,
14'b00011100010011,
14'b00110000011000,
14'b00111000111111,
14'b00101110111111,
14'b00000010101011,
14'b00001110110100,
14'b01000111111010,
14'b00100111010011,
14'b01000111000001,
14'b00111100111111,
14'b00110001011011,
14'b00101010111011,
14'b00000001101001,
14'b00011111100100,
14'b01000001001010,
14'b00001001111111,
14'b00010001101001,
14'b00010101011111,
14'b00100111000110,
14'b00001010100010,
14'b00100101111111,
14'b00011001011001,
14'b00000110110001,
14'b00110101111000,
14'b00001100001100,
14'b00011001110110,
14'b01000001101110,
14'b00001101000100,
14'b00011110110011,
14'b00110000100111,
14'b00001010001001,
14'b00111000000110,
14'b01000000110110,
14'b00111000010000,
14'b00110111001100,
14'b00001101001001,
14'b00111110101101,
14'b01000010001001,
14'b00000100000000,
14'b01000011110010,
14'b00100011101011,
14'b00100101110111,
14'b00101001000100,
14'b00001011111110,
14'b00111100011010,
14'b01000001100001,
14'b00000111001110,
14'b00101110010110,
14'b00000000101110,
14'b00111000110100,
14'b00100011101101,
14'b00011111000100,
14'b00100000110100,
14'b00001100000111,
14'b00011100000000,
14'b00110010101111,
14'b00101010111101,
14'b00100100111010,
14'b00000100100000,
14'b00010011010001,
14'b00010111101001,
14'b00111111110110,
14'b00110110001111,
14'b00110001110110,
14'b00011001111000,
14'b00111011011111,
14'b00000010001101,
14'b01000010111100,
14'b00011110011010,
14'b00011101101100,
14'b00111011010101,
14'b00110100100111,
14'b00111101101011,
14'b00101001110110,
14'b00000111010110,
14'b00011010011111,
14'b00101111010101,
14'b00100100000011,
14'b00010111000001,
14'b00000100000100,
14'b00110100001011,
14'b00110101100001,
14'b00011100110001,
14'b00010100010000,
14'b00000111101111,
14'b00011100100110,
14'b00000100110100,
14'b00110100010000,
14'b00010011111011,
14'b00100101011100,
14'b00101000000001,
14'b01000100100100,
14'b00011101011100,
14'b00011101011110,
14'b00101111011000,
14'b00010010011111,
14'b00001101000101,
14'b00101100010110,
14'b00010100000011,
14'b00000100001100,
14'b00011011010101,
14'b00011010111111,
14'b00000010100111,
14'b01000000011000,
14'b01000001111111,
14'b00101111001110,
14'b00101010111001,
14'b00101111111010,
14'b00000110010111,
14'b00111100101111,
14'b00100100001101,
14'b00100000001000,
14'b00011110011011,
14'b01000111000000,
14'b00100101011011,
14'b00001000111001,
14'b00011000011001,
14'b00011111111100,
14'b00110001101100,
14'b00001001000010,
14'b00101010001111,
14'b00101110110100,
14'b00000010011001,
14'b00010110101110,
14'b00111010010000,
14'b00110000011010,
14'b00111101111111,
14'b00000111111110,
14'b00011010110100,
14'b00101001100111,
14'b00010011110001,
14'b01000110111001,
14'b01000000110101,
14'b00100101000010,
14'b00010101100111,
14'b00010111111100,
14'b00010110010011,
14'b00010101111100,
14'b00010101111001,
14'b00000010011011,
14'b00001101111001,
14'b00100110111101,
14'b00011001101101,
14'b00100100111000,
14'b00011100100001,
14'b00011111000010,
14'b00010110110000,
14'b00101101010100,
14'b01000001111011,
14'b01000010110110,
14'b00001100110011,
14'b00001101110110,
14'b00101011000011,
14'b00101010011110,
14'b01000001001111,
14'b01000101011000,
14'b00011101010001,
14'b00001101111011,
14'b00000011000111,
14'b00110101011001,
14'b00101101101101,
14'b00111111000001,
14'b00011010011010,
14'b01000011010100,
14'b01000010110000,
14'b00101111010000,
14'b00110011011101,
14'b00111011011011,
14'b00101100010100,
14'b00011110010010,
14'b00000110000000,
14'b01000111111110,
14'b00011101010100,
14'b00111110010010,
14'b00111010011000,
14'b00110100011001,
14'b00011000100111,
14'b01000111010110,
14'b00010110100000,
14'b00001111000110,
14'b00110000101010,
14'b00011001010101,
14'b01000010000010,
14'b00001011001101,
14'b00111010101010,
14'b00111101110111,
14'b00011010001101,
14'b00010110001000,
14'b00111011010011,
14'b00100000100100,
14'b00100101111101,
14'b00001001011111,
14'b00010010000100,
14'b00011011000111,
14'b00000101000011,
14'b00100100011110,
14'b00111111000100,
14'b01000001001001,
14'b00000001110100,
14'b00101011010111,
14'b01000000010010,
14'b00011001100101,
14'b00111000101110,
14'b00000000000101,
14'b00101010100011,
14'b00011110111110,
14'b00010000111111,
14'b00111010100111,
14'b00111110100100,
14'b00010000001011,
14'b00101110111010,
14'b01000110110011,
14'b00101011011111,
14'b00000110111101,
14'b00011001101010,
14'b00111010101111,
14'b00100101100001,
14'b00000010001010,
14'b00111110010101,
14'b00000100011101,
14'b00100100100001,
14'b00010101110111,
14'b00000000000110,
14'b00111000011100,
14'b00001110010000,
14'b00110100011101,
14'b00111011011000,
14'b00111000100011,
14'b00010000100110,
14'b00110001101110,
14'b00111011101101,
14'b00111111001101,
14'b00101110010001,
14'b01000010010000,
14'b00010110111110,
14'b00111010001001,
14'b00001000000001,
14'b00111001000011,
14'b00100100110101,
14'b00010111001010,
14'b00001101111000,
14'b00001111001010,
14'b01000101000011,
14'b00000100011010,
14'b00100111011111,
14'b00000111111011,
14'b00111100011000,
14'b00110011010001,
14'b01000111111111,
14'b00110000011100,
14'b00000111101100,
14'b00000000100001,
14'b00010101101000,
14'b00101001111000,
14'b00011101111010,
14'b00000100010000,
14'b01000000100100,
14'b00001111011111,
14'b01000101010000,
14'b01000010100011,
14'b00110010010000,
14'b00101111010100,
14'b00000101111110,
14'b00010101110011,
14'b00111010010100,
14'b00011101011111,
14'b00111011001011,
14'b00010100011011,
14'b00010100011101,
14'b00010011100110,
14'b00101111001011,
14'b01000100011110,
14'b00011011101010,
14'b00111010100010,
14'b00111110000000,
14'b00001111010101,
14'b00011110100001,
14'b00001111000100,
14'b00001010110000,
14'b00111000101111,
14'b01000001011001,
14'b00011010000010,
14'b00010101000000,
14'b00011001001101,
14'b00001011101001,
14'b00001010101011,
14'b00010111001111,
14'b00111110011001,
14'b00000110000111,
14'b00010001010011,
14'b00001000011001,
14'b00000001100000,
14'b00011000001101,
14'b00111010010101,
14'b00010001101101,
14'b01000111111011,
14'b00100110011111,
14'b00100111111100,
14'b00100100110111,
14'b00011110110001,
14'b00010000010000,
14'b00001111010000,
14'b00010101010011,
14'b00110011000011,
14'b00010010100101,
14'b00110111011110,
14'b01000001110101,
14'b00101110001100,
14'b00010010011001,
14'b00111110101010,
14'b00100010111001,
14'b00100011010110,
14'b00100011010100,
14'b00111110110110,
14'b00110001010011,
14'b00110001001010,
14'b00100101010100,
14'b01000111101010,
14'b00011111110110,
14'b00001101001101,
14'b00100110011011,
14'b00110010000110,
14'b00110010011011,
14'b00000100011111,
14'b00100010110111,
14'b00010110011110,
14'b00000101101100,
14'b00111110101011,
14'b00111110110100,
14'b00100011010101,
14'b00010001100000,
14'b00101110011001,
14'b00111011001110,
14'b00111101101001,
14'b00110011011100,
14'b00111001010100,
14'b00001101100010,
14'b00100100110001,
14'b00111100001110,
14'b00001110000011,
14'b00001011111010,
14'b00001111010111,
14'b00100100010001,
14'b01000100011111,
14'b00010011100111,
14'b00001110000100,
14'b00110001011010,
14'b00101010000101,
14'b00000110011011,
14'b01000111001001,
14'b00011100101011,
14'b00000111110111,
14'b00011011110100,
14'b00001100000010,
14'b00011000101011,
14'b00001011001100,
14'b00100110001010,
14'b00111001001100,
14'b01000001101011,
14'b00000001011001,
14'b00011001001111,
14'b00111011011110,
14'b00100101001100,
14'b00011100111111,
14'b00001010010011,
14'b00000100001101,
14'b00000001101101,
14'b00111100000100,
14'b00011010100001,
14'b00001110000010,
14'b00100111011110,
14'b01000101100010,
14'b00100010110100,
14'b00110000000011,
14'b00101001011010,
14'b00110011011000,
14'b00111101111011,
14'b00010011110101,
14'b00100011001111,
14'b00010001010101,
14'b00110010010101,
14'b00111100111001,
14'b00010111011100,
14'b01000110100010,
14'b00100011111010,
14'b00101010110011,
14'b00011010101010,
14'b00100101101111,
14'b00010101110110,
14'b00111110010100,
14'b00000111000001,
14'b00111010100011,
14'b00011110110000,
14'b00101100110000,
14'b00001011000001,
14'b00101001001000,
14'b00100001101011,
14'b00010111010111,
14'b00011111010001,
14'b00010111111111,
14'b00010111101101,
14'b00111000001100,
14'b00100011010011,
14'b00111101011101,
14'b00100000101110,
14'b00010011011000,
14'b00111110100101,
14'b00111110110111,
14'b00000011101101,
14'b00001100011110,
14'b00000000011110,
14'b00110001010101,
14'b00111111011100,
14'b00100111010010,
14'b00000101001001,
14'b00001111110000,
14'b00011111111111,
14'b00001110000110,
14'b00000101010110,
14'b00011100110010,
14'b00101111001111,
14'b00010010100100,
14'b01000011001001,
14'b00100001101111,
14'b00110010011001,
14'b00011000001011,
14'b00001001100010,
14'b00111000010100,
14'b00101110111101,
14'b00110110010010,
14'b00110011010011,
14'b01000110001010,
14'b00010010001010,
14'b00100111001111,
14'b01000010010011,
14'b00110001000011,
14'b00101100010111,
14'b00100011011010,
14'b00101110100011,
14'b00000101011101,
14'b00111011010000,
14'b00111100010000,
14'b01000110000101,
14'b00100101110001,
14'b00010101100011,
14'b00100000001110,
14'b00101100100000,
14'b00110101110011,
14'b00100111111101,
14'b00111110011100,
14'b00001100100110,
14'b00111101001110,
14'b00111110001101,
14'b00010100011100,
14'b00101010001110,
14'b00110100110100,
14'b01000011010000,
14'b00000010111000,
14'b00010000001001,
14'b00100100010110,
14'b00001110011011,
14'b00110111100011,
14'b01000010111011,
14'b00111100110110,
14'b00001011110111,
14'b01000111011001,
14'b00110001011111,
14'b00111010011011,
14'b00111011111110,
14'b00101010111111,
14'b00000001010100,
14'b00001111011101,
14'b00010010101110,
14'b00010001111101,
14'b00011011010010,
14'b00010011000110,
14'b00110101110110,
14'b00110101110001,
14'b01000011010101,
14'b00111010111101,
14'b00110001111101,
14'b00101110101011,
14'b00110111001010,
14'b00011011011100,
14'b00110110001000,
14'b00110111110010,
14'b01000101100011,
14'b00100001001101,
14'b00011101100010,
14'b01000000001000,
14'b01000010001101,
14'b00000001111111,
14'b01000110110010,
14'b00011110010111,
14'b01000001001101,
14'b01000100111010,
14'b01000011100011,
14'b00010011011111,
14'b00010010010000,
14'b00100000011101,
14'b00110110100111,
14'b00001111000111,
14'b00010000000010,
14'b00000110100111,
14'b00001101011100,
14'b00110010000101,
14'b00101111011010,
14'b00010100101101,
14'b00001000100101,
14'b00000010000100,
14'b00111001111001,
14'b01000010100001,
14'b01000101010010,
14'b00001101000001,
14'b00101110101111,
14'b00011110000011,
14'b00011011110101,
14'b00101110101000,
14'b00010100110001,
14'b01000100110000,
14'b01001000000000,
14'b00101000011111,
14'b00010111110011,
14'b00000110110010,
14'b00001101011011,
14'b00010111101000,
14'b00101000100101,
14'b00101100011111,
14'b01000111000011,
14'b00010000011011,
14'b00111010110100,
14'b00000010100010,
14'b00000010110101,
14'b00000110111100,
14'b01000101000110,
14'b00101001101100,
14'b00100010010000,
14'b00101000111011,
14'b00101101001110,
14'b01000010110010,
14'b00010011110100,
14'b00101011111110,
14'b00110011001111,
14'b00111111010110,
14'b00110100110111,
14'b00101010001001,
14'b01000110110100,
14'b00011101111110,
14'b00110001000001,
14'b00001100100011,
14'b00100111011001,
14'b00111100001011,
14'b00011101010010,
14'b00010001110101,
14'b00001100101111,
14'b00110010001001,
14'b01000100001010,
14'b00010101010110,
14'b00000011111011,
14'b00101000101011,
14'b00101000111101,
14'b00000001000101,
14'b00111111100011,
14'b00000010011101,
14'b00001100100000,
14'b00011001110100,
14'b00100110111111,
14'b00011010010001,
14'b01000010010111,
14'b00101011110001,
14'b00001111100001,
14'b00110010110110,
14'b00010000010101,
14'b00000001101000,
14'b00010110101000,
14'b00110111011100,
14'b00100100110100,
14'b00001001011101,
14'b00010101100100,
14'b00111110001001,
14'b00111100001100,
14'b00010011000111,
14'b00111000000101,
14'b00001000011010,
14'b00001011001010,
14'b00111011000100,
14'b00001110101011,
14'b01000100001001,
14'b00100001111001,
14'b00111001001101,
14'b01000111100011,
14'b00111101010001,
14'b00000000011111,
14'b00100000011110,
14'b00000110111000,
14'b00100110101111,
14'b00111101011000,
14'b00110011011110,
14'b00101110010010,
14'b00100011010000,
14'b00000011000001,
14'b00101101010111,
14'b00001000110011,
14'b00001011011111,
14'b00000110000011,
14'b00010111100111,
14'b00101111101001,
14'b01000010011000,
14'b00100001000100,
14'b00100111000100,
14'b00110001010000,
14'b00001000100111,
14'b00011100111101,
14'b00010001110000,
14'b00100101110101,
14'b00110101110010,
14'b00001000101001,
14'b00010100110111,
14'b00111001011000,
14'b00110010110100,
14'b00100100000111,
14'b00010011111101,
14'b00011010110110,
14'b00011100000101,
14'b00110101100010,
14'b00110010100001,
14'b00001101100000,
14'b00100101001110,
14'b00110011101001,
14'b00111101110010,
14'b00010100110101,
14'b00101000010100,
14'b00000100101101,
14'b00010110001110,
14'b00010101101110,
14'b01000000110000,
14'b00000101011100,
14'b00011101111001,
14'b00110001010110,
14'b00010011001101,
14'b00101110011100,
14'b00011001101001,
14'b00011000101000,
14'b00111001011001,
14'b00111011111001,
14'b01000011001000,
14'b00110100000110,
14'b01000100011101,
14'b00001010010111,
14'b00111001001001,
14'b00101100100011,
14'b01000110010011,
14'b01000111001111,
14'b01000101010111,
14'b00011110111101,
14'b00111110100001,
14'b00110100001000,
14'b00010000011000,
14'b00101101101010,
14'b00010001011101,
14'b00001000011100,
14'b00100001111011,
14'b00100110010001,
14'b00101001001111,
14'b00000011111010,
14'b00010010011011,
14'b00100100001001,
14'b00001101110001,
14'b00101001110011,
14'b00010111100011,
14'b00110111110110,
14'b00101010001010,
14'b01000010011010,
14'b00101110011011,
14'b00010100010100,
14'b00001010010000,
14'b00001111010010,
14'b00001101110010,
14'b00100101000111,
14'b00011100101110,
14'b01000110100101,
14'b00100110110010,
14'b00001101111111,
14'b00011000011110,
14'b00010010101001,
14'b00011100101010,
14'b00101000110100,
14'b01000101100001,
14'b00101111000110,
14'b00010000000011,
14'b00001110001001,
14'b00100000011000,
14'b00000110011010,
14'b00010111011010,
14'b00110001011001,
14'b00001110001010,
14'b00110011001001,
14'b00111111011111,
14'b00100110100100,
14'b00000101001101,
14'b00101110101100,
14'b01000010000111,
14'b00010110011101,
14'b00010011000010,
14'b00110000110010,
14'b00110100011100,
14'b00001100110000,
14'b00000101101000,
14'b00101100001110,
14'b00111000001101,
14'b01000100000010,
14'b01000000110100,
14'b00111101110000,
14'b00101100000001};