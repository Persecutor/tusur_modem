(* ram_style = "block" *) logic [11:0] map_i [0:1023] = {
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010100000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010100000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010100000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010100000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010101000,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b101010101010,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b101010101010,
12'b000000000000,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b010101010101,
12'b101010101010,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b010101010100,
12'b101010101000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010100000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010100000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010100000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b010101010000,
12'b101010100000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b010101000000,
12'b101010000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b010100000000,
12'b101000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b010000000000,
12'b100000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000};
