logic [23:0] sig_pr [0:2047] = {
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000000111111111111,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000001000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b111111111111000000000000,
24'b000000001100000000000101,
24'b000000000001000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000101,
24'b000000000001000000000000,
24'b000000001101000000000111,
24'b000000000000000000000001,
24'b000000001011000000000101,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000101,
24'b000000000001000000000000,
24'b000000001100000000000110,
24'b000000000000111111111111,
24'b000000001101000000000110,
24'b111111111111000000000001,
24'b000000001100000000000100,
24'b000000000001000000000000,
24'b000000001101000000000110,
24'b000000000000000000000001,
24'b000000001100000000000101,
24'b000000000000000000000001,
24'b000000001100000000000101,
24'b000000000001000000000001,
24'b000000001100000000000101,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b111111111111000000000000,
24'b000000001100000000000101,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001101000000000101,
24'b111111111111000000000000,
24'b000000001101000000000100,
24'b111111111111000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000001000000000001,
24'b000000001101000000000101,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000001,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000001,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000001000000000000,
24'b000000001110000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000000,
24'b000000001110000000000100,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001101000000000100,
24'b000000000000111111111111,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001110000000000011,
24'b000000000000111111111111,
24'b000000001111000000000100,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000001000000000001,
24'b000000001110000000000100,
24'b000000000001000000000000,
24'b000000001111000000000100,
24'b000000000000000000000001,
24'b000000001110000000000100,
24'b111111111111000000000000,
24'b000000001110000000000011,
24'b000000000000000000000000,
24'b000000001110000000000010,
24'b000000000000111111111111,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000010000000000000011,
24'b000000000000000000000000,
24'b000000001111000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000001000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000001111000000000011,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000001000000000000,
24'b000000010000000000000011,
24'b000000000000000000000000,
24'b000000010001000000000010,
24'b000000000001000000000000,
24'b000000010001000000000011,
24'b000000000001000000000001,
24'b000000010000000000000011,
24'b000000000000000000000000,
24'b000000010000000000000011,
24'b111111111111000000000000,
24'b000000010001000000000010,
24'b000000000000000000000000,
24'b000000010000000000000010,
24'b000000000000000000000000,
24'b000000010001000000000010,
24'b000000000000000000000000,
24'b000000010001000000000010,
24'b000000000000000000000000,
24'b000000010000000000000001,
24'b000000000000111111111111,
24'b000000010010000000000010,
24'b000000000000000000000001,
24'b000000010001000000000010,
24'b111111111111000000000000,
24'b000000010001000000000001,
24'b000000000000000000000000,
24'b000000010010000000000001,
24'b000000000000000000000000,
24'b000000010010000000000010,
24'b000000000000000000000000,
24'b000000010010000000000001,
24'b000000000000000000000001,
24'b000000010001000000000001,
24'b111111111111000000000000,
24'b000000010010000000000000,
24'b000000000000000000000001,
24'b000000010001000000000001,
24'b000000000000000000000000,
24'b000000010010000000000001,
24'b111111111111000000000000,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000001,
24'b000000000000000000000000,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000000,
24'b000000000000000000000001,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000000,
24'b000000000001000000000001,
24'b000000010010000000000000,
24'b000000000000000000000000,
24'b000000010011000000000000,
24'b000000000001000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100000000000000,
24'b000000000000000000000000,
24'b000000010100111111111111,
24'b000000000001000000000000,
24'b000000010100000000000000,
24'b111111111111000000000000,
24'b000000010100111111111111,
24'b000000000000000000000000,
24'b000000010100111111111111,
24'b000000000001000000000000,
24'b000000010100000000000000,
24'b111111111111000000000000,
24'b000000010100111111111111,
24'b000000000001111111111111,
24'b000000010101000000000000,
24'b000000000000111111111111,
24'b000000010110111111111111,
24'b000000000000000000000000,
24'b000000010110111111111111,
24'b111111111111000000000000,
24'b000000010101111111111110,
24'b000000000001111111111111,
24'b000000010110111111111111,
24'b000000000000000000000000,
24'b000000010110111111111110,
24'b000000000000000000000000,
24'b000000010111111111111111,
24'b111111111111000000000000,
24'b000000010111111111111111,
24'b000000000000000000000000,
24'b000000010111111111111111,
24'b111111111111000000000000,
24'b000000010111111111111110,
24'b111111111111111111111111,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011001111111111110,
24'b000000000000000000000001,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011000111111111110,
24'b000000000000000000000000,
24'b000000011001111111111101,
24'b000000000000000000000000,
24'b000000011001111111111101,
24'b000000000000000000000000,
24'b000000011010111111111101,
24'b000000000000000000000000,
24'b000000011001111111111101,
24'b000000000001111111111111,
24'b000000011010111111111110,
24'b000000000000000000000000,
24'b000000011011111111111101,
24'b111111111111000000000000,
24'b000000011011111111111100,
24'b000000000000000000000001,
24'b000000011010111111111101,
24'b000000000000111111111111,
24'b000000011100111111111101,
24'b000000000000000000000000,
24'b000000011100111111111101,
24'b000000000000000000000000,
24'b000000011100111111111101,
24'b111111111111000000000000,
24'b000000011101111111111100,
24'b000000000000000000000000,
24'b000000011101111111111101,
24'b111111111111000000000000,
24'b000000011110111111111100,
24'b000000000000000000000000,
24'b000000011110111111111101,
24'b111111111111000000000000,
24'b000000011111111111111100,
24'b111111111111000000000000,
24'b000000011111111111111011,
24'b000000000000000000000000,
24'b000000100000111111111011,
24'b000000000000000000000001,
24'b000000100000111111111100,
24'b000000000000000000000000,
24'b000000100001111111111011,
24'b000000000000000000000000,
24'b000000100001111111111011,
24'b000000000000000000000000,
24'b000000100010111111111011,
24'b000000000000000000000001,
24'b000000100010111111111011,
24'b000000000000000000000000,
24'b000000100011111111111010,
24'b000000000000000000000000,
24'b000000100100111111111011,
24'b111111111111000000000000,
24'b000000100101111111111010,
24'b111111111111000000000000,
24'b000000100110111111111001,
24'b000000000000000000000001,
24'b000000100110111111111010,
24'b000000000000000000000000,
24'b000000100111111111111010,
24'b000000000000000000000000,
24'b000000101001111111111010,
24'b000000000000000000000001,
24'b000000101001111111111010,
24'b111111111111000000000000,
24'b000000101010111111111001,
24'b111111111111000000000000,
24'b000000101010111111111000,
24'b000000000000111111111111,
24'b000000101100111111111001,
24'b111111111111111111111111,
24'b000000101110111111111000,
24'b000000000000000000000000,
24'b000000101111111111111000,
24'b111111111111000000000000,
24'b000000110001111111111000,
24'b000000000000000000000001,
24'b000000110001111111110111,
24'b000000000000000000000000,
24'b000000110011111111110111,
24'b000000000000000000000000,
24'b000000110101111111110110,
24'b000000000000000000000000,
24'b000000110111111111110110,
24'b000000000000000000000001,
24'b000000111000111111110110,
24'b000000000000000000000000,
24'b000000111011111111110110,
24'b000000000000000000000001,
24'b000000111101111111110101,
24'b000000000000000000000000,
24'b000000111110111111110101,
24'b000000000000111111111111,
24'b000001000011111111110100,
24'b000000000000000000000000,
24'b000001000110111111110100,
24'b000000000000000000000000,
24'b000001001001111111110011,
24'b000000000000000000000000,
24'b000001001100111111110010,
24'b000000000000000000000000,
24'b000001010001111111110000,
24'b000000000001000000000000,
24'b000001010101111111101111,
24'b000000000000111111111111,
24'b000001011011111111101110,
24'b111111111111000000000000,
24'b000001100001111111101010,
24'b000000000000000000000000,
24'b000001101001111111100111,
24'b111111111111000000000000,
24'b000001110000111111100010,
24'b000000000000000000000000,
24'b000001111010111111011011,
24'b000000000001000000000001,
24'b000010000100111111010001,
24'b000000000000000000000000,
24'b000010010000111111000000,
24'b000000000000000000000000,
24'b000010011100111110100000,
24'b000000000000000000000000,
24'b000010011010111101010110,
24'b000000000000000000000000,
24'b111111010111110111111011,
24'b001011010110110100101010,
24'b010100001011000010010110,
24'b001011010110001011010110,
24'b000110111001010000001110,
24'b110100101010001011010110,
24'b000001000111111000000011,
24'b001011010110001011010110,
24'b110101000100001110010001,
24'b110100101001110100101001,
24'b010000000010110111100000,
24'b001011010101001011010101,
24'b000100101001001110011010,
24'b110100101001001011010110,
24'b000000110111111000010101,
24'b001011010101001011010101,
24'b111101111000010000100110,
24'b110100101010001011010110,
24'b111010000010000010100110,
24'b110100101010001011010110,
24'b101110011101110101000000,
24'b001011010101110100101010,
24'b001001000001001111000111,
24'b110100101010001011010110,
24'b111011110101000010111011,
24'b110100101001001011010111,
24'b101110010011111110000010,
24'b110100101010110100101010,
24'b000111101111111000110001,
24'b110100101010001011010110,
24'b111001010001101010110000,
24'b001011010110001011010110,
24'b101001010001111010100110,
24'b001011010110110100101010,
24'b110111101101000010110011,
24'b001011010110110100101001,
24'b111101100110010010100111,
24'b110100101011110100101010,
24'b000011011000000100100010,
24'b110100101001110100101010,
24'b010001011101111111000111,
24'b110100101010001011010101,
24'b000000101100111010000011,
24'b110100101010001011010101,
24'b110000010011101101100100,
24'b001011010101110100101010,
24'b000000000010000111001010,
24'b110100101011110100101010,
24'b001111010010111000101011,
24'b110100101010001011010111,
24'b111000001110101000100010,
24'b001011010110110100101010,
24'b010000100001110110110010,
24'b001011010110001011010110,
24'b000011100010111100011000,
24'b001011010110001011010111,
24'b111110001100000001101001,
24'b001011010110001011010110,
24'b111000100110001110011101,
24'b110100101001001011010110,
24'b101010010001110101110010,
24'b001011010110110100101010,
24'b111001110011001011101001,
24'b110100101001110100101011,
24'b000001100000110100100001,
24'b001011010110110100101010,
24'b010000100000001010111111,
24'b110100101010001011010110,
24'b000000100001110100001100,
24'b001011010110001011010101,
24'b110001100011001010111010,
24'b110100101010110100101010,
24'b001001011011110100100001,
24'b001011010110001011010110,
24'b110011010000001100010100,
24'b110100101010110100101010,
24'b001010011001111101100011,
24'b110100101010001011010110,
24'b110100010111101110101001,
24'b001011010110110100101010,
24'b001100101011000101111101,
24'b110100101011001011010110,
24'b111111000101101110001010,
24'b001011010110001011010110,
24'b110111111011111100100000,
24'b001011010110001011010111,
24'b101000101011001010011110,
24'b110100101010110100101010,
24'b110111001010110000111111,
24'b001011010110110100101010,
24'b111100111001111110110011,
24'b001011010111110100101010,
24'b000010011010001100110101,
24'b110100101010110100101001,
24'b010000001010110100010100,
24'b001011010110001011010111,
24'b111110110100001001110110,
24'b110100101010001011010110,
24'b101101100011110001100001,
24'b001011010110110100101010,
24'b111011011011000000000001,
24'b001011010110110100101010,
24'b000001101101001111011000,
24'b110100101010110100101010,
24'b001110011100111110111111,
24'b110100101011001011010101,
24'b110100101111101111010001,
24'b001011010110110100101001,
24'b000010110111000101110111,
24'b110100101010110100101001,
24'b010010001001101101001001,
24'b001011010111001011010101,
24'b000001111010111001100111,
24'b001011010110001011010110,
24'b110010011111111110001101,
24'b001011010111110100101010,
24'b001001101011000010101000,
24'b001011010110001011011000,
24'b110001111110001110011001,
24'b110100101010110100101010,
24'b000000110101110011101110,
24'b001011010110110100101010,
24'b010000010110000000000001,
24'b001011010110001011010110,
24'b111111110110000110001100,
24'b001011010111001011010110,
24'b101111001010010100011100,
24'b110100101010110100101010,
24'b111101101110000100100111,
24'b110100101010110100101010,
24'b000101000100111100011010,
24'b110100101001110100101010,
24'b010100001100101100100011,
24'b001011010110001011010110,
24'b000101011010111010101010,
24'b001011010111001011010111,
24'b111111001010000000001011,
24'b001011010111001011010110,
24'b111000110100000101101000,
24'b001011010110001011010111,
24'b101001101001010011011101,
24'b110100101010110100101010,
24'b110111111011000010100110,
24'b110100101010110100101011,
24'b111101000011110010110010,
24'b001011010111110100101010,
24'b000000111100001001101001,
24'b110100101010110100101010,
24'b000101011111110001100011,
24'b001011010110110100101010,
24'b010001110110111111101110,
24'b001011010101001011010110,
24'b111000101111001101101000,
24'b110100101010110100101001,
24'b001101111101110100001111,
24'b001011010110001011010110,
24'b110101010000000010011000,
24'b001011010110110100101001,
24'b000010101100010001100000,
24'b110100101010110100101011,
24'b001001110101000000110001,
24'b110100101010110100101010,
24'b011001001110110000000011,
24'b001011010110001011010110,
24'b001011000110111111001011,
24'b001011010110001011010110,
24'b000110001100001101010011,
24'b110100101001001011010110,
24'b000010110001110011110111,
24'b001011010101001011010110,
24'b111111011111000001101010,
24'b001011010101001011010111,
24'b111011000011001111100001,
24'b110100101010001011010111,
24'b101110000000110110010100,
24'b001011010101110100101010,
24'b111111110110000100110110,
24'b001011010110110100101010,
24'b010001101011010100110011,
24'b110100101010001011010110,
24'b000100101000000110000101,
24'b110100101010001011010110,
24'b000000001101111111001101,
24'b110100101010001011010101,
24'b111100111101110001111011,
24'b001011010110001011010101,
24'b111001100100001011001001,
24'b110100101011001011010110,
24'b110100110000111100011110,
24'b110100101001001011010110,
24'b100110111001101100010111,
24'b001011010110110100101010,
24'b110111010000111011000001,
24'b001011010110110100101011,
24'b000101110110000010000101,
24'b001011010110001011010110,
24'b101100010010010000011001,
24'b110100101011110100101010,
24'b111000111000111111011101,
24'b110100101010110100101010,
24'b111110100000101110100110,
24'b001011010110110100101001,
24'b001010100101111101100101,
24'b001011010101001011010110,
24'b101111101100001011011100,
24'b110100101010110100101010,
24'b111011001110110001100001,
24'b001011010110110100101010,
24'b111111001000111110000001,
24'b001011010110110100101010,
24'b000010010111000011111001,
24'b001011010101110100101010,
24'b000110100001010000101011,
24'b110100101010110100101001,
24'b010010101101110111110011,
24'b001011010110001011010110,
24'b111001100111001101011010,
24'b110100101001110100101010,
24'b001111001100110101111101,
24'b001011010101001011010110,
24'b110111111001001011111011,
24'b110100101010110100101010,
24'b001110010001110100011110,
24'b001011010110001011010110,
24'b110111100110001010000001,
24'b110100101010110100101010,
24'b001111000101110001000011,
24'b001011010110001011010110,
24'b111111110010111101100100,
24'b001011010110001011010111,
24'b101111011111000010100000,
24'b001011010110110100101010,
24'b111110001100000111101000,
24'b001011010111110100101010,
24'b000101100011010101010010,
24'b110100101010110100101010,
24'b010100100011000100001010,
24'b110100101010001011010110,
24'b000101011000110011100011,
24'b001011010110001011010101,
24'b111101111000000011010011,
24'b001011010110001011010111,
24'b101110111101010011011010,
24'b110100101010110100101010,
24'b111110111101000100010110,
24'b110100101010110100101001,
24'b001101110011111100100000,
24'b110100101010001011010110,
24'b110101000110101100110011,
24'b001011010110110100101010,
24'b000011111111111010110100,
24'b001011010110110100101010,
24'b010100001010111111111001,
24'b001011010110001011010110,
24'b000101100110000011111000,
24'b001011010110001011010101,
24'b111110110010001000110000,
24'b001011010110001011010111,
24'b110001010110010110001111,
24'b110100101010110100101010,
24'b001001101101000100111100,
24'b110100101001001011010110,
24'b110011101010110011110111,
24'b001011010110110100101010,
24'b001010101000000010001110,
24'b001011010110001011010110,
24'b110100000011001001011100,
24'b001011010110110100101010,
24'b001010101111011000010110,
24'b110100101010001011010110,
24'b110011111010001000101001,
24'b110100101010110100101010,
24'b001010001110111010100001,
24'b001011010110001011010110,
24'b110010010111010100100100,
24'b110100101010110100101010,
24'b000001001110001000101101,
24'b110100101010110100101010,
24'b010000110100000100110001,
24'b110100101010001011010110,
24'b000000011111000001111000,
24'b110100101010001011010111,
24'b110000001001111111000000,
24'b110100101011110100101010,
24'b111111110001111011000110,
24'b110100101010110100101001,
24'b001110101110101111010010,
24'b001011010110001011010101,
24'b110111001001001001011100,
24'b110100101010110100101010,
24'b001110011010111011011011,
24'b110100101010001011010110,
24'b111111000101101011110111,
24'b001011010110001011010110,
24'b101110111100111010111011,
24'b001011010111110100101011,
24'b111110010111000010010001,
24'b001011010110110100101010,
24'b001100101101010000010011,
24'b110100101001001011010110,
24'b110011011010111000110101,
24'b001011010110110100101010,
24'b000001010001010000111001,
24'b110100101010110100101011,
24'b001111000110000011100111,
24'b110100101010001011010111,
24'b110101101101111101010111,
24'b110100101011110100101010,
24'b000011110011110000100001,
24'b001011010101110100101001,
24'b010010010100001010000010,
24'b110100101010001011010101,
24'b111010110010111011101010,
24'b110100101001110100101011,
24'b010010100011101011110111,
24'b001011010110001011010110,
24'b000100110101111010110111,
24'b001011010110001011010110,
24'b111101110101000010011010,
24'b001011010110001011010110,
24'b101111001100010001100010,
24'b110100101011110100101010,
24'b111111010101000010011111,
24'b110100101010110100101010,
24'b001110001100111011001010,
24'b110100101010001011010110,
24'b110101011101101101000100,
24'b001011010110110100101010,
24'b000100001100000100010010,
24'b110100101011110100101010,
24'b010011111001101011110101,
24'b001011010111001011010101,
24'b000011111000111000010011,
24'b001011010110001011010110,
24'b110100000110111100100100,
24'b001011010110110100101010,
24'b000100101001111111110110,
24'b001011010110110100101010,
24'b010101101011000011101101,
24'b001011010110001011010111,
24'b000111111011001111000101,
24'b110100101010001011010110,
24'b000010100110110011111011,
24'b001011010110001011010110,
24'b111101010011111111011101,
24'b001011010111001011010110,
24'b101111101101000011101111,
24'b001011010110110100101010,
24'b000000111111001000001111,
24'b001011010110110100101010,
24'b010010000000010100100101,
24'b110100101011001011010101,
24'b000011000001111011100111,
24'b001011010110001011010110,
24'b110100110101010001010001,
24'b110100101010110100101011,
24'b001101011101111010000100,
24'b001011010110001011010101,
24'b111000011000010000100001,
24'b110100101010110100101010,
24'b010001100110111001110101,
24'b001011010101001011010110,
24'b000101001010010000110000,
24'b110100101010001011010101,
24'b111111110001111010110000,
24'b001011010110001011010110,
24'b110011111010010011010010,
24'b110100101010110100101011,
24'b001110111100000110001100,
24'b110100101010001011010110,
24'b000011100100000000000010,
24'b110100101010001011010110,
24'b111111101101110011000101,
24'b001011010110001011010110,
24'b111100011100001011111110,
24'b110100101010001011010101,
24'b111000000010110110101001,
24'b001011010111001011010110,
24'b101010110011001111010000,
24'b110100101010110100101010,
24'b111100000100000001010010,
24'b110100101010110100101010,
24'b001100001100110011011100,
24'b001011010110001011010110,
24'b110101101101001100111010,
24'b110100101010110100101010,
24'b001110010101111110111101,
24'b110100101010001011010111,
24'b000001010110110000101011,
24'b001011010110001011010110,
24'b111011010010001000101011,
24'b110100101010001011010110,
24'b101110010110110010001110,
24'b001011010110110100101010,
24'b000111000100001000011100,
24'b110100101011001011010110,
24'b110001010011101111111111,
24'b001011010111110100101010,
24'b001000100000111100111011,
24'b001011010110001011010110,
24'b110010000111000010001011,
24'b001011010110110100101001,
24'b001000110101000111100001,
24'b001011010110001011010110,
24'b110001011011010100110010,
24'b110100101010110100101010,
24'b000000110101111101000101,
24'b001011010110110100101010,
24'b010001010100010101001101,
24'b110100101010001011010110,
24'b000010111010001000011110,
24'b110100101010001011010110,
24'b111100000010000011111101,
24'b110100101011001011010110,
24'b101101110111000000100011,
24'b110100101010110100101010,
24'b111111000001111101000010,
24'b110100101010110100101001,
24'b010000010100111000000101,
24'b110100101010001011010111,
24'b000010100111101001111110,
24'b001011010110001011010110,
24'b111101001101111001011010,
24'b001011010110001011010111,
24'b110111101101000000100111,
24'b001011010110001011010111,
24'b101001101100001110000010,
24'b110100101011110100101010,
24'b111010010001110100110110,
24'b001011010110110100101010,
24'b001001100110000011011010,
24'b001011010110001011010101,
24'b110001111111010011001011,
24'b110100101001110100101010,
24'b001000010011000011011110,
24'b110100101010001011010110,
24'b110001010000110100111010,
24'b001011010110110100101001,
24'b000111011000001101111111,
24'b110100101010001011010111,
24'b101111001101111111110000,
24'b110100101010110100101010,
24'b111101011111110001001110,
24'b001011010110110100101010,
24'b001011100100001000111000,
24'b110100101010001011010110,
24'b110010010111110001011100,
24'b001011010110110100101010,
24'b000000101111000000001011,
24'b001011010110110100101010,
24'b010000001010001110101011,
24'b110100101001001011010110,
24'b111111111110110101111011,
24'b001011010110001011010101,
24'b110000100011000100111100,
24'b001011010111110100101010,
24'b000111100101010101011100,
24'b110100101001001011010110,
24'b101111011110000111100000,
24'b110100101001110100101001,
24'b111101000000000010010100,
24'b110100101010110100101010,
24'b000011110101111110000110,
24'b110100101010110100101010,
24'b010010011000111000101111,
24'b110100101011001011010110,
24'b000010001000101010010110,
24'b001011010110001011010110,
24'b110011000001111001011001,
24'b001011010110110100101010,
24'b001010111011111111100111,
24'b001011010110001011010110,
24'b110101000101000101101011,
24'b001011010101110100101010,
24'b001101011101010100000110,
24'b110100101010001011010110,
24'b111111111011000011111010,
24'b110100101001001011010110,
24'b111000110101110100111010,
24'b001011010110001011010110,
24'b101001110001001100111101,
24'b110100101010110100101010,
24'b111000101001110111001111,
24'b001011010111110100101010,
24'b111111100001001111101011,
24'b110100101001110100101010,
24'b001100110101000001101000,
24'b110100101010001011010110,
24'b110100001100110011111011,
24'b001011010110110100101010,
24'b001001101100001101110001,
24'b110100101001001011010101,
24'b110001010011000000111110,
24'b110100101010110100101011,
24'b111111100011111010100011,
24'b110100101001110100101100,
24'b001101111001101100010101,
24'b001011010111001011010110,
24'b110101111110111101000100,
24'b001011010110110100101010,
24'b001100111100001101010100,
24'b110100101010001011010101,
24'b111101010100111101001001,
24'b110100101010001011010110,
24'b101100101010101100011111,
24'b001011010110110100101010,
24'b111010111001111010110001,
24'b001011010111110100101011,
24'b000001011011000001010111,
24'b001011010111110100101010,
24'b001110100011001110011110,
24'b110100101010001011010110,
24'b110101111001110101100111,
24'b001011010111110100101011,
24'b001011100010001010110001,
24'b110100101010001011010110,
24'b110100000011110001101100,
24'b001011010111110100101010,
24'b001001101111111110001111,
24'b001011010110001011010110,
24'b110001000101000011001100,
24'b001011010111110100101010,
24'b111110010011001000010010,
24'b001011010110110100101010,
24'b000100111110010101010001,
24'b110100101011110100101011,
24'b010011100001111101001100,
24'b001011010110001011010110,
24'b000011111100010100101010,
24'b110100101010001011010110,
24'b111011111011000110010000,
24'b110100101010001011010110,
24'b101100010010111000100000,
24'b001011010110110100101010,
24'b111010101110010010100110,
24'b110100101010110100101010,
24'b000001001001000110100101,
24'b110100101011110100101010,
24'b001101110001000010010000,
24'b110100101010001011010101,
24'b110011100110111110100001,
24'b110100101010110100101010,
24'b000000001110111001100100,
24'b110100101010110100101010,
24'b000110100110101011100100,
24'b001011010111110100101010,
24'b010100110111111011001101,
24'b001011010111001011010111,
24'b000100011011000010110000,
24'b001011010101001011010101,
24'b110101010111010000101110,
24'b110100101010110100101010,
24'b001101111010111000111100,
24'b001011010101001011010110,
24'b111111000000001111100111,
24'b110100101010001011010110,
24'b101111000010111001100100,
24'b001011010111110100101010,
24'b111110100101010001111101,
24'b110100101010110100101010,
24'b001100111111000100000011,
24'b110100101010001011010110,
24'b110011110001110110100001,
24'b001011010110110100101010,
24'b000001110000010000100001,
24'b110100101010110100101010,
24'b001111110011000011011011,
24'b110100101010001011010110,
24'b110110110000110110100100,
24'b001011010110110100101010,
24'b000101011111010001011110,
24'b110100101010110100101001,
24'b010101101110000110010010,
24'b110100101011001011010110,
24'b000111011101000011000000,
24'b110100101010001011010110,
24'b000001101110000000110110,
24'b110100101001001011010110,
24'b111100000101111111000010,
24'b110100101010001011010101,
24'b101110001000111101010011,
24'b110100101010110100101010,
24'b111111000010111011011000,
24'b110100101010110100101011,
24'b001111100010111000111110,
24'b110100101010001011010110,
24'b111111111101110101001100,
24'b110100101010001011010111,
24'b110000110110101001000101,
24'b001011010110110100101010,
24'b001000000101000001111000,
24'b110100101010001011010110,
24'b110000000101101011000100,
24'b001011010110110100101001,
24'b111101100100111010001101,
24'b001011010110110100101010,
24'b000100000111001001000001,
24'b110100101001110100101010,
24'b010001100011110000111101,
24'b001011010111001011010110,
24'b111001011001000110101110,
24'b110100101010110100101010,
24'b001111111011101110001101,
24'b001011010110001011010110,
24'b111001110111111011011111,
24'b001011010110110100101010,
24'b010010100111000010001001,
24'b001011010110001011010110,
24'b000110001010010000011000,
24'b110100101010001011010111,
24'b000001101111111111100010,
24'b110100101010001011010110,
24'b111110010101101110111100,
24'b001011010111001011010101,
24'b111010110001111110010110,
24'b001011010110001011010110,
24'b110101101011001101000001,
24'b110100101010001011010110,
24'b100111010100110100111010,
24'b001011010110110100101010,
24'b110110001111001010110001,
24'b110100101010110100101010,
24'b111100001111110010101101,
24'b001011010110110100101010,
24'b000001111000000001011111,
24'b001011010111110100101010,
24'b001111101010010001000101,
24'b110100101010001011010110,
24'b111110010101000000110011,
24'b110100101010001011010110,
24'b101100111110110000100111,
24'b001011010110110100101010,
24'b111010101010000000011010,
24'b001011010110110100101100,
24'b000000100100001111101001,
24'b110100101010110100101001,
24'b001100110000111000100010,
24'b001011010110001011010110,
24'b110001111011010000101000,
24'b110100101010110100101011,
24'b111101011100000011001101,
24'b110100101010110100101010,
24'b000001010101111100100010,
24'b110100101010110100101010,
24'b000100011000101110010101,
24'b001011010110110100101010,
24'b000111101010111111010000,
24'b001011010110110100101010,
24'b001100011011010000000001,
24'b110100101001110100101001,
24'b011010000101000001000010,
24'b110100101010001011010110,
24'b000110110100110101101111,
24'b000000000000000000000000,
24'b010000001111110110111100,
24'b001011010110001011010100,
24'b001000001011001010011101,
24'b110100101010001011010101,
24'b000100011110110010101100,
24'b001011010110001011010110,
24'b000001001110000001111011,
24'b001011010101001011010110,
24'b111101001000010010001000,
24'b110100101010001011010110,
24'b110001001010000010111000,
24'b110100101001110100101010,
24'b001010101100110100110101,
24'b001011010110001011010111,
24'b110110000000001110110000,
24'b110100101010110100101010,
24'b001111011110000010011100,
24'b110100101010001011010110,
24'b000011010101111101011111,
24'b110100101011001011010110,
24'b111110110101111000001001,
24'b110100101010001011010110,
24'b111010011000101010000011,
24'b001011010110001011010110,
24'b101110011011111001110101,
24'b001011010110110100101011,
24'b001000110011000001111000,
24'b001011010111001011010110,
24'b111100000010010001100100,
24'b110100101001001011010101,
24'b110101001111000011001011,
24'b110100101010001011010101,
24'b100110000010111101010111,
24'b110100101010110100101010,
24'b110100001100110111100000,
24'b110100101010110100101010,
24'b111001000110101001000101,
24'b001011010111110100101001,
24'b111100011011111001000101,
24'b001011010110110100101001,
24'b111111011100000111011011,
24'b110100101011110100101010,
24'b000011010000101101100111,
24'b001011010110110100101010,
24'b001110101000111001101101,
24'b001011010110001011010110,
24'b110011100010111101111111,
24'b001011010110110100101001,
24'b111111001010000001010010,
24'b001011010110110100101001,
24'b000011100100000100110011,
24'b001011010110110100101010,
24'b001000001110001001110100,
24'b001011010110110100101010,
24'b010100110100011000000011,
24'b110100101001001011010101,
24'b111100011000001000110001,
24'b110100101001110100101011,
24'b010011010111000001101110,
24'b110100101010001011010101,
24'b000100010110110100011101,
24'b001011010110001011010110,
24'b110101100010001101010011,
24'b110100101010110100101010,
24'b001101010111111000010010,
24'b001011010110001011010101,
24'b110111000011010001101001,
24'b110100101001110100101010,
24'b001101110000000101100111,
24'b110100101010001011010110,
24'b110110011010000001100110,
24'b110100101011110100101010,
24'b000110000010111110101001,
24'b110100101010110100101011,
24'b010110111011111011100011,
24'b110100101011001011010110,
24'b001001011011110111001100,
24'b110100101010001011010101,
24'b000100110101101001111101,
24'b001011010111001011010110,
24'b000001100011111011011000,
24'b001011010110001011010110,
24'b111110010011001100010001,
24'b110100101010001011010110,
24'b111001110101111100110111,
24'b110100101010001011010110,
24'b101100100101101101011000,
24'b001011010110110100101010,
24'b111110000010111110000100,
24'b001011010110110100101011,
24'b001111000100001111000101,
24'b110100101010001011010110,
24'b000000000100000001001100,
24'b110100101010001011010110,
24'b110001111000111011100011,
24'b110100101010110100101010,
24'b001011000100110101101110,
24'b110100101011001011010101,
24'b111100101011100111001100,
24'b001011010110001011010110,
24'b101101001100110110011000,
24'b001011010111110100101011,
24'b111101001111111101101011,
24'b001011010110110100101011,
24'b001100011010001100000001,
24'b110100101011001011010110,
24'b110100111100111010111010,
24'b110100101010110100101010,
24'b001100001011101001100000,
24'b001011010110001011010110,
24'b111100101000110110110110,
24'b001011010110001011010101,
24'b101011111011111011100000,
24'b001011010110110100101010,
24'b111001101100111111001010,
24'b001011010110110100101010,
24'b111110101011000011101101,
24'b001011010110110100101001,
24'b000010101000010000110100,
24'b110100101010110100101010,
24'b000111010111111110111111,
24'b110100101011110100101011,
24'b010100000011101101001011,
24'b001011010110001011010110,
24'b111011100010111010001111,
24'b001011010111110100101010,
24'b010001110110111110110000,
24'b001011010110001011010110,
24'b111011101001000010010001,
24'b001011010110110100101011,
24'b010100001101000110101000,
24'b001011010111001011010110,
24'b000111010110010010111101,
24'b110100101010001011010110,
24'b000001101000111010000001,
24'b001011010110001011010111,
24'b110101100100001111110010,
24'b110100101010110100101010,
24'b010000100000111000101100,
24'b001011010111001011010110,
24'b000101000101001111011001,
24'b110100101010001011010110,
24'b000001010010111001001000,
24'b001011010110001011010101,
24'b111110010000010001010011,
24'b110100101001001011010111,
24'b111010011000000011001010,
24'b110100101001001011010110,
24'b101110110010110101011101,
24'b001011010110110100101010,
24'b001001010100001111011111,
24'b110100101010001011010110,
24'b111100000111000011001111,
24'b110100101010001011010111,
24'b101110100101111110010100,
24'b110100101011110100101010,
24'b000111111111111001000001,
24'b110100101010001011010110,
24'b111001011111101010111100,
24'b001011010110001011010110,
24'b101001011111111010110001,
24'b001011010110110100101001,
24'b110111111011000010111011,
24'b001011010101110100101001,
24'b111101110100010010101101,
24'b110100101010110100101011,
24'b000011100100000100100101,
24'b110100101010110100101010,
24'b010001101010111111001010,
24'b110100101010001011010110,
24'b000000110111111010000101,
24'b110100101010001011010110,
24'b110000011101101101100100,
24'b001011010110110100101010,
24'b000000001100000111001010,
24'b110100101011110100101010,
24'b001111011010111000101001,
24'b110100101010001011010101,
24'b111000011000101000100001,
24'b001011010110110100101011,
24'b010000101000110110101111,
24'b001011010110001011010101,
24'b000011101010111100010100,
24'b001011010110001011010110,
24'b111110010101000001100100,
24'b001011010110001011010110,
24'b111000101110001110011000,
24'b110100101010001011010110,
24'b101010011000110101101101,
24'b001011010110110100101001,
24'b111001111010001011100011,
24'b110100101010110100101010,
24'b000001100111110100011100,
24'b001011010110110100101001,
24'b010000101000001010111000,
24'b110100101010001011010110,
24'b000000101000110100000101,
24'b001011010110001011010101,
24'b110001101011001010110010,
24'b110100101010110100101010,
24'b001001100001110100011001,
24'b001011010110001011010101,
24'b110011010111001100001100,
24'b110100101010110100101010,
24'b001010011111111101011010,
24'b110100101010001011010101,
24'b110100011111101110100000,
24'b001011010110110100101011,
24'b001100110001000101110100,
24'b110100101011001011010110,
24'b111111001100101110000001,
24'b001011010110001011010110,
24'b111000000000111100010111,
24'b001011010110001011010110,
24'b101000110001001010010100,
24'b110100101001110100101010,
24'b110111010000110000110101,
24'b001011010110110100101010,
24'b111100111111111110101001,
24'b001011010110110100101011,
24'b000010011111001100101010,
24'b110100101010110100101010,
24'b010000001110110100001001,
24'b001011010110001011010110,
24'b111110111010001001101011,
24'b110100101001001011010110,
24'b101101101000110001010101,
24'b001011010111110100101010,
24'b111011100000111111110111,
24'b001011010110110100101010,
24'b000001110001001111001101,
24'b110100101010110100101010,
24'b001110100010111110110100,
24'b110100101010001011010110,
24'b110100110101101111000100,
24'b001011010110110100101011,
24'b000010111011000101101011,
24'b110100101011110100101010,
24'b010010001101101100111110,
24'b001011010110001011010110,
24'b000001111101111001011001,
24'b001011010111001011010110,
24'b110010100010111110000001,
24'b001011010110110100101010,
24'b001001101110000010011100,
24'b001011010101001011010110,
24'b110010000011001110001100,
24'b110100101010110100101001,
24'b000000111011110011100000,
24'b001011010110110100101011,
24'b010000011010111111110101,
24'b001011010110001011010110,
24'b111111111010000110000000,
24'b001011010101001011010101,
24'b101111001111010100001110,
24'b110100101010110100101011,
24'b111101110010000100011001,
24'b110100101010110100101010,
24'b000101000111111100001101,
24'b110100101010110100101001,
24'b010100010000101100010110,
24'b001011010110001011010110,
24'b000101011110111010011101,
24'b001011010110001011010111,
24'b111111001110111111111110,
24'b001011010110001011010111,
24'b111000110111000101011010,
24'b001011010110001011010110,
24'b101001101101010011001111,
24'b110100101010110100101010,
24'b110111111111000010011000,
24'b110100101010110100101010,
24'b111101001000110010100101,
24'b001011010101110100101011,
24'b000001000000001001011001,
24'b110100101011110100101010,
24'b000101100010110001010101,
24'b001011010110110100101010,
24'b010001111001111111100000,
24'b001011010111001011010110,
24'b111000110010001101011011,
24'b110100101010110100101010,
24'b001110000000110100000001,
24'b001011010110001011010110,
24'b110101010011000010001011,
24'b001011010101110100101010,
24'b000010101110010001010001,
24'b110100101001110100101010,
24'b001001111000000000100011,
24'b110100101001110100101010,
24'b011001010001101111110100,
24'b001011010110001011010110,
24'b001011001010111110111011,
24'b001011010110001011010111,
24'b000110001111001101000100,
24'b110100101010001011010111,
24'b000010110010110011101000,
24'b001011010110001011010101,
24'b111111100001000001011100,
24'b001011010110001011010101,
24'b111011000111001111010011,
24'b110100101010001011010101,
24'b101110000100110110000101,
24'b001011010110110100101010,
24'b111111111001000100101000,
24'b001011010101110100101001,
24'b010001101111010100100100,
24'b110100101010001011010111,
24'b000100101011000101110110,
24'b110100101011001011010101,
24'b000000010001111110111110,
24'b110100101010001011010110,
24'b111101000000110001101100,
24'b001011010110001011010110,
24'b111001100110001010111010,
24'b110100101010001011010101,
24'b110100110011111100001110,
24'b110100101010001011010110,
24'b100110111100101100001000,
24'b001011010111110100101010,
24'b110111010010111010110010,
24'b001011010110110100101001,
24'b000101111001000001110110,
24'b001011010111001011010101,
24'b101100010110010000001011,
24'b110100101001110100101010,
24'b111000111101111111001101,
24'b110100101010110100101011,
24'b111110100100101110010111,
24'b001011010110110100101010,
24'b001010101000111101010101,
24'b001011010110001011010110,
24'b101111101111001011001101,
24'b110100101010110100101010,
24'b111011010000110001010001,
24'b001011010111110100101010,
24'b111111001100111101110010,
24'b001011010110110100101010,
24'b000010011011000011101001,
24'b001011010110110100101011,
24'b000110100100010000011100,
24'b110100101001110100101011,
24'b010010101110110111100100,
24'b001011010110001011010101,
24'b111001101001001101001010,
24'b110100101010110100101001,
24'b001111001111110101101101,
24'b001011010110001011010110,
24'b110111111100001011101101,
24'b110100101010110100101010,
24'b001110010100110100001111,
24'b001011010110001011010110,
24'b110111101001001001110010,
24'b110100101010110100101010,
24'b001111001000110000110100,
24'b001011010101001011010110,
24'b111111110101111101010100,
24'b001011010110001011010111,
24'b101111100010000010001111,
24'b001011010110110100101011,
24'b111110001110000111011001,
24'b001011010110110100101010,
24'b000101100101010101000010,
24'b110100101010110100101010,
24'b010100100111000011111010,
24'b110100101010001011010110,
24'b000101011011110011010010,
24'b001011010110001011010110,
24'b111101111010000011000011,
24'b001011010110001011010110,
24'b101111000000010011001010,
24'b110100101010110100101010,
24'b111111000001000100000110,
24'b110100101010110100101001,
24'b001101110110111100001111,
24'b110100101010001011010110,
24'b110101001001101100100001,
24'b001011010110110100101011,
24'b000100000001111010100100,
24'b001011010110110100101010,
24'b010100001101111111101001,
24'b001011010101001011010110,
24'b000101101001000011100111,
24'b001011010110001011010110,
24'b111110110011001000011111,
24'b001011010110001011010110,
24'b110001011000010101111110,
24'b110100101001110100101010,
24'b001001110000000100101010,
24'b110100101010001011010101,
24'b110011101101110011100111,
24'b001011010101110100101010,
24'b001010101011000001111101,
24'b001011010110001011010111,
24'b110100000110001001001010,
24'b001011010110110100101010,
24'b001010110001011000000101,
24'b110100101010001011010110,
24'b110011111110001000010111,
24'b110100101010110100101010,
24'b001010010001111010001111,
24'b001011010110001011010110,
24'b110010011010010100010010,
24'b110100101010110100101010,
24'b000001010010001000011011,
24'b110100101011110100101010,
24'b010000110110000100011111,
24'b110100101011001011010110,
24'b000000100001000001100110,
24'b110100101011001011010110,
24'b110000001101111110101111,
24'b110100101010110100101010,
24'b111111110101111010110101,
24'b110100101010110100101010,
24'b001110110001101111000001,
24'b001011010101001011010110,
24'b110111001100001001001001,
24'b110100101010110100101010,
24'b001110011101111011000111,
24'b110100101011001011010111,
24'b111111000111101011100101,
24'b001011010111001011010101,
24'b101110111111111010101010,
24'b001011010110110100101010,
24'b111110011011000001111111,
24'b001011010110110100101010,
24'b001100110000001111111111,
24'b110100101010001011010110,
24'b110011011100111000100011,
24'b001011010110110100101010,
24'b000001010100010000100110,
24'b110100101010110100101010,
24'b001111001001000011010011,
24'b110100101011001011010101,
24'b110101110010111101000101,
24'b110100101010110100101011,
24'b000011110110110000001101,
24'b001011010110110100101010,
24'b010010010110001001101111,
24'b110100101010001011010101,
24'b111010110100111011010111,
24'b110100101010110100101010,
24'b010010100110101011100100,
24'b001011010110001011010110,
24'b000100111000111010100100,
24'b001011010110001011010101,
24'b111101111010000010000110,
24'b001011010110001011010111,
24'b101111001111010001001111,
24'b110100101010110100101010,
24'b111111011000000010001011,
24'b110100101001110100101010,
24'b001110010000111010110101,
24'b110100101010001011010110,
24'b110101100001101100110000,
24'b001011010110110100101010,
24'b000100010000000011111110,
24'b110100101010110100101010,
24'b010011111101101011100000,
24'b001011010110001011010110,
24'b000011111100110111111101,
24'b001011010110001011010111,
24'b110100000111111100010000,
24'b001011010110110100101001,
24'b000100101100111111100000,
24'b001011010101110100101001,
24'b010101101111000011010111,
24'b001011010110001011010111,
24'b000111111111001110101111,
24'b110100101010001011010110,
24'b000010101010110011100110,
24'b001011010110001011010111,
24'b111101010111111111000111,
24'b001011010101001011010110,
24'b101111110001000011011000,
24'b001011010111110100101011,
24'b000001000011000111111001,
24'b001011010110110100101010,
24'b010010000011010100001110,
24'b110100101010001011010101,
24'b000011000101111011001111,
24'b001011010110001011010110,
24'b110100111000010000111010,
24'b110100101001110100101001,
24'b001101100011111001101011,
24'b001011010111001011010110,
24'b111000011100010000001010,
24'b110100101011110100101010,
24'b010001101010111001011101,
24'b001011010111001011010110,
24'b000101001110010000011001,
24'b110100101010001011010101,
24'b111111110101111010011000,
24'b001011010110001011010110,
24'b110011111101010010111010,
24'b110100101011110100101001,
24'b001111000010000101110100,
24'b110100101010001011010111,
24'b000011101000111111101010,
24'b110100101010001011010110,
24'b111111110010110010101101,
24'b001011010110001011010110,
24'b111100100010001011100100,
24'b110100101010001011010111,
24'b111000000101110110010001,
24'b001011010110001011010110,
24'b101010110111001110110110,
24'b110100101010110100101010,
24'b111100001000000000111000,
24'b110100101010110100101010,
24'b001100010001110011000011,
24'b001011010101001011010111,
24'b110101110001001100100000,
24'b110100101010110100101010,
24'b001110011000111110100011,
24'b110100101001001011010110,
24'b000001011011110000001111,
24'b001011010110001011010101,
24'b111011010111001000010000,
24'b110100101010001011010101,
24'b101110011100110001110010,
24'b001011010110110100101010,
24'b000111001010001000000000,
24'b110100101010001011010110,
24'b110001011001101111100010,
24'b001011010110110100101010,
24'b001000100110111100011110,
24'b001011010110001011010111,
24'b110010001100000001101110,
24'b001011010110110100101010,
24'b001000111010000111000100,
24'b001011010110001011010110,
24'b110001100000010100010100,
24'b110100101001110100101010,
24'b000000111010111100100101,
24'b001011010111110100101001,
24'b010001011010010100101111,
24'b110100101010001011010101,
24'b000011000000001000000000,
24'b110100101010001011010110,
24'b111100001000000011011110,
24'b110100101010001011010110,
24'b101101111110000000000011,
24'b110100101010110100101010,
24'b111111001000111100100001,
24'b110100101010110100101010,
24'b010000011001110111100100,
24'b110100101010001011010110,
24'b000010101110101001011101,
24'b001011010110001011010110,
24'b111101010100111000111000,
24'b001011010110001011010110,
24'b110111110101000000000101,
24'b001011010101001011010110,
24'b101001110101001101011111,
24'b110100101001110100101010,
24'b111010011001110100010000,
24'b001011010111110100101010,
24'b001001101111000010110110,
24'b001011010111001011010110,
24'b110010000111010010100111,
24'b110100101001110100101011,
24'b001000011011000010111001,
24'b110100101001001011010111,
24'b110001011000110100010100,
24'b001011010110110100101010,
24'b000111100000001101011000,
24'b110100101010001011011000,
24'b101111010100111111001001,
24'b110100101010110100101001,
24'b111101101001110000100111,
24'b001011010110110100101010,
24'b001011101100001000010000,
24'b110100101011001011010110,
24'b110010100000110000110010,
24'b001011010111110100101010,
24'b000000111000111111100010,
24'b001011010110110100101001,
24'b010000010101001110000000,
24'b110100101010001011010111,
24'b000000001000110101001111,
24'b001011010111001011010101,
24'b110000101110000100010000,
24'b001011010110110100101010,
24'b000111110000010100101111,
24'b110100101010001011010110,
24'b101111101010000110110010,
24'b110100101001110100101010,
24'b111101001010000001100101,
24'b110100101010110100101010,
24'b000100000001111101010110,
24'b110100101010110100101010,
24'b010010100101111000000000,
24'b110100101001001011010110,
24'b000010010100101001100011,
24'b001011010110001011010110,
24'b110011001111111000100101,
24'b001011010110110100101010,
24'b001011001001111110110010,
24'b001011010111001011010110,
24'b110101010011000100110101,
24'b001011010110110100101010,
24'b001101101011010011001111,
24'b110100101010001011010110,
24'b000000001010000011000001,
24'b110100101010001011010110,
24'b111001000110110100000000,
24'b001011010110001011010110,
24'b101010000010001100000001,
24'b110100101010110100101010,
24'b111000111011110110010010,
24'b001011010110110100101010,
24'b111111110100001110101011,
24'b110100101001110100101010,
24'b001101001001000000100111,
24'b110100101010001011010110,
24'b110100100010110010111000,
24'b001011010110110100101010,
24'b001010000010001100101100,
24'b110100101010001011010110,
24'b110001101001111111110111,
24'b110100101010110100101010,
24'b111111111011111001011001,
24'b110100101010110100101010,
24'b001110010101101011001001,
24'b001011010110001011010110,
24'b110110011011111011110101,
24'b001011010110110100101001,
24'b001101011101001100000010,
24'b110100101010001011010111,
24'b111101110101111011110011,
24'b110100101010001011010110,
24'b101101010000101011000111,
24'b001011010110110100101011,
24'b111011100001111001010101,
24'b001011010111110100101010,
24'b000010001000111111110111,
24'b001011010110110100101010,
24'b001111010110001100111000,
24'b110100101011001011010110,
24'b110110110011110011111110,
24'b001011010110110100101010,
24'b001100101001001001000100,
24'b110100101010001011010111,
24'b110101011000101111111110,
24'b001011010110110100101010,
24'b001011100011111100100100,
24'b001011010110001011010110,
24'b110100000000000001111100,
24'b001011010110110100101011,
24'b000110011011001010110010,
24'b000000000001000000000000,
24'b000010001100000100101100,
24'b000000000000000000000000,
24'b000001011100000011001000,
24'b000000000000000000000000,
24'b000001000110000010011000,
24'b000000000000000000000000,
24'b000000111010000001111011,
24'b000000000000000000000000,
24'b000000110001000001100111,
24'b000000000000000000000000,
24'b000000101011000001011000,
24'b000000000000000000000000,
24'b000000100111000001001101,
24'b000000000001000000000000,
24'b000000100011000001000110,
24'b000000000000000000000000,
24'b000000100000000000111111,
24'b000000000000000000000000,
24'b000000011101000000111010,
24'b000000000000000000000000,
24'b000000011011000000110101,
24'b000000000000000000000000,
24'b000000011001000000110001,
24'b000000000000111111111111,
24'b000000011000000000101110,
24'b000000000000000000000000,
24'b000000010111000000101011,
24'b000000000001000000000000,
24'b000000010101000000101001,
24'b000000000000000000000001,
24'b000000010100000000100111,
24'b000000000000000000000001,
24'b000000010010000000100110,
24'b111111111111000000000000,
24'b000000010001000000100011,
24'b000000000000111111111111,
24'b000000010010000000100010,
24'b111111111111000000000000,
24'b000000010000000000100000,
24'b000000000000000000000000,
24'b000000010000000000011111,
24'b000000000000000000000001,
24'b000000001110000000011110,
24'b000000000000000000000000,
24'b000000001110000000011101,
24'b000000000000000000000000,
24'b000000001110000000011100,
24'b000000000000000000000000,
24'b000000001101000000011011,
24'b000000000000000000000000,
24'b000000001100000000011010,
24'b000000000001000000000000,
24'b000000001100000000011010,
24'b000000000000111111111111,
24'b000000001100000000011010,
24'b111111111111000000000000,
24'b000000001100000000011001,
24'b111111111111000000000000,
24'b000000001100000000011000,
24'b000000000000000000000001,
24'b000000001010000000010111,
24'b000000000000111111111111,
24'b000000001011000000010111,
24'b000000000001000000000000,
24'b000000001011000000010111,
24'b111111111111000000000000,
24'b000000001010000000010110,
24'b000000000000000000000000,
24'b000000001011000000010101,
24'b000000000000000000000000,
24'b000000001010000000010101,
24'b000000000000000000000000,
24'b000000001010000000010100,
24'b000000000000000000000000,
24'b000000001001000000010101,
24'b000000000000000000000000,
24'b000000001010000000010100,
24'b000000000000000000000000,
24'b000000001010000000010100,
24'b000000000000000000000001,
24'b000000001001000000010100,
24'b000000000000000000000000,
24'b000000001001000000010011,
24'b000000000000000000000000,
24'b000000001001000000010011,
24'b000000000000000000000000,
24'b000000001001000000010011,
24'b111111111111000000000000,
24'b000000001001000000010010,
24'b000000000000000000000000,
24'b000000001001000000010010,
24'b000000000000000000000000,
24'b000000001000000000010010,
24'b000000000000000000000000,
24'b000000001000000000010001,
24'b000000000000000000000000,
24'b000000001001000000010001,
24'b000000000000000000000001,
24'b000000000111000000010001,
24'b000000000000000000000000,
24'b000000000111000000010001,
24'b000000000000111111111111,
24'b000000001000000000010001,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000001,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000000111000000010000,
24'b000000000000000000000000,
24'b000000001000000000010000,
24'b000000000000000000000000,
24'b000000000111000000001111,
24'b000000000000111111111111,
24'b000000000111000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b111111111111000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000000111000000001111,
24'b000000000000000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000000,
24'b000000001000000000001111,
24'b000000000000000000000001,
24'b000000000111000000001110,
24'b000000000000000000000000,
24'b000000000111000000001110,
24'b000000000000000000000000,
24'b000000000111000000001110,
24'b000000000000000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000000111000000001110,
24'b111111111111000000000000,
24'b000000001000000000001110,
24'b000000000000000000000000,
24'b000000000111000000001101,
24'b000000000000000000000000,
24'b000000001000000000001101,
24'b000000000000000000000000,
24'b000000000111000000001101,
24'b111111111111111111111111,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000001000000000001101,
24'b111111111111000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000001000000000001101,
24'b111111111111000000000001,
24'b000000000111000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000001,
24'b000000000111000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000000111000000001100,
24'b000000000001000000000000,
24'b000000001000000000001101,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000000000000000,
24'b000000000111000000001100,
24'b111111111111000000000000,
24'b000000000111000000001100,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b111111111111000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000000111000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001100,
24'b000000000000111111111111,
24'b000000001000000000001011,
24'b000000000001000000000001,
24'b000000001000000000001100,
24'b111111111111000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000111111111111,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000000000000000,
24'b000000001000000000001011,
24'b000000000000111111111111,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000111111111111,
24'b000000001000000000001010,
24'b000000000000111111111111,
24'b000000001001000000001010,
24'b000000000001000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000001000000000000,
24'b000000001001000000001011,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000001,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001000000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000000,
24'b000000001001000000001010,
24'b000000000000000000000001,
24'b000000001000000000001010,
24'b111111111111000000000000,
24'b000000001001000000001010,
24'b111111111111000000000000,
24'b000000001000000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b111111111111000000000000,
24'b000000001010000000001001,
24'b000000000000000000000001,
24'b000000001000000000001001,
24'b000000000000111111111111,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001010000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000001000000000001,
24'b000000001001000000001001,
24'b000000000000000000000000,
24'b000000001001000000001001,
24'b000000000000111111111111,
24'b000000001001000000001001,
24'b111111111111111111111111,
24'b000000001001000000001001,
24'b111111111111111111111111,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b111111111111000000000001,
24'b000000001001000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000001,
24'b000000001010000000001000,
24'b111111111111000000000000,
24'b000000001010000000000111,
24'b000000000001000000000000,
24'b000000001010000000001000,
24'b111111111111000000000000,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000001,
24'b000000001001000000000111,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b000000000001000000000001,
24'b000000001001000000001000,
24'b111111111111111111111111,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001010000000001000,
24'b000000000000111111111111,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001011000000001000,
24'b111111111111000000000000,
24'b000000001010000000000110,
24'b000000000001000000000000,
24'b000000001011000000001000,
24'b111111111111000000000001,
24'b000000001010000000000111,
24'b000000000000111111111111,
24'b000000001011000000000111,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b111111111111000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b000000000000111111111111,
24'b000000001011000000000111,
24'b000000000000000000000000,
24'b000000001011000000000110,
24'b000000000001000000000000,
24'b000000001011000000000111,
24'b000000000000000000000001,
24'b000000001011000000000111,
24'b000000000000000000000000,
24'b000000001011000000000111,
24'b111111111111000000000000,
24'b000000001011000000000110,
24'b000000000000000000000000,
24'b000000001010000000000111,
24'b111111111111111111111111,
24'b000000001100000000000110,
24'b000000000000000000000000,
24'b000000001100000000000110,
24'b000000000001000000000001,
24'b000000001010000000000111};