logic [1:0] map_p [0:1023] = {
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b00,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b11,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00,
2'b00}