(* ram_style = "block" *) logic [11:0] map_p [0:1023] = {
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b000000000000,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111111,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111111100,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111110000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111111000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b111100000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b110000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000,
12'b000000000000};