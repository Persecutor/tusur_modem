logic [23:0] sig_pr [0:2047] = {
24'b111111111111000000000000,
24'b000000001010111111111000,
24'b000000000000000000000000,
24'b000000001010111111111000,
24'b000000000000111111111111,
24'b000000001011111111110111,
24'b000000000011000000000000,
24'b000000001011111111111011,
24'b000000000000000000000000,
24'b000000001011111111111010,
24'b111111111111000000000000,
24'b000000001100111111111001,
24'b111111111111000000000001,
24'b000000001011111111111001,
24'b111111111111000000000001,
24'b000000001010111111111000,
24'b000000000001111111111111,
24'b000000001011111111111001,
24'b000000000000111111111111,
24'b000000001100111111111010,
24'b111111111110000000000001,
24'b000000001011111111111000,
24'b000000000000000000000001,
24'b000000001011111111111001,
24'b111111111111000000000000,
24'b000000001010111111111000,
24'b111111111110000000000000,
24'b000000001011111111110110,
24'b000000000000000000000000,
24'b000000001011111111111000,
24'b000000000000000000000000,
24'b000000001011111111111000,
24'b111111111111000000000000,
24'b000000001010111111110111,
24'b000000000001111111111111,
24'b000000001011111111111000,
24'b111111111111111111111111,
24'b000000001100111111110111,
24'b000000000001111111111111,
24'b000000001100111111111000,
24'b000000000001111111111111,
24'b000000001101111111111000,
24'b000000000001000000000000,
24'b000000001101111111111000,
24'b000000000001000000000000,
24'b000000001100111111111001,
24'b111111111111000000000000,
24'b000000001101111111110111,
24'b000000000001111111111111,
24'b000000001101111111111001,
24'b000000000001000000000001,
24'b000000001100111111111001,
24'b111111111111111111111111,
24'b000000001101111111111000,
24'b000000000000000000000000,
24'b000000001101111111111001,
24'b111111111111000000000000,
24'b000000001101111111111000,
24'b111111111111000000000000,
24'b000000001110111111110111,
24'b000000000000000000000000,
24'b000000001110111111111001,
24'b111111111110000000000000,
24'b000000001110111111110110,
24'b000000000000000000000001,
24'b000000001101111111110111,
24'b000000000001111111111111,
24'b000000001110111111111000,
24'b111111111111000000000001,
24'b000000001110111111110110,
24'b000000000000000000000000,
24'b000000001101111111110111,
24'b000000000000111111111111,
24'b000000001110111111110111,
24'b000000000000111111111111,
24'b000000001111111111110111,
24'b000000000010000000000001,
24'b000000001110111111111000,
24'b000000000000000000000000,
24'b000000001111111111111000,
24'b000000000000111111111111,
24'b000000010000111111111000,
24'b000000000000000000000001,
24'b000000001110111111111000,
24'b000000000000111111111111,
24'b000000010000111111111000,
24'b000000000000000000000000,
24'b000000010000111111111000,
24'b111111111110000000000000,
24'b000000010000111111110111,
24'b111111111111000000000001,
24'b000000001111111111110110,
24'b000000000000000000000000,
24'b000000010001111111110111,
24'b111111111111000000000001,
24'b000000001111111111110110,
24'b111111111111000000000001,
24'b000000010000111111110101,
24'b000000000000000000000001,
24'b000000001111111111110101,
24'b000000000001000000000000,
24'b000000010000111111110110,
24'b000000000001000000000000,
24'b000000010000111111110111,
24'b111111111111111111111111,
24'b000000010010111111110101,
24'b000000000001000000000000,
24'b000000010010111111111000,
24'b111111111111000000000001,
24'b000000010000111111110110,
24'b000000000000111111111111,
24'b000000010010111111110110,
24'b000000000000000000000000,
24'b000000010001111111110111,
24'b000000000000111111111111,
24'b000000010011111111110111,
24'b111111111111000000000000,
24'b000000010010111111110110,
24'b000000000000111111111111,
24'b000000010100111111110110,
24'b000000000000000000000001,
24'b000000010010111111110111,
24'b111111111110111111111111,
24'b000000010011111111110100,
24'b000000000001111111111111,
24'b000000010100111111110101,
24'b000000000001000000000000,
24'b000000010100111111110110,
24'b000000000000111111111111,
24'b000000010110111111110110,
24'b000000000000000000000001,
24'b000000010101111111110110,
24'b111111111111000000000001,
24'b000000010100111111110101,
24'b000000000000000000000000,
24'b000000010110111111110101,
24'b111111111111000000000001,
24'b000000010101111111110101,
24'b000000000000000000000000,
24'b000000010101111111110101,
24'b000000000000000000000000,
24'b000000010110111111110101,
24'b111111111111000000000000,
24'b000000010111111111110100,
24'b000000000000000000000000,
24'b000000010111111111110100,
24'b000000000000000000000001,
24'b000000010101111111110101,
24'b000000000000111111111110,
24'b000000011000111111110100,
24'b000000000010000000000000,
24'b000000011000111111110111,
24'b111111111101111111111111,
24'b000000011010111111110100,
24'b111111111111000000000000,
24'b000000011010111111110100,
24'b111111111111000000000001,
24'b000000011001111111110010,
24'b000000000001000000000000,
24'b000000011010111111110101,
24'b000000000000000000000000,
24'b000000011011111111110100,
24'b111111111111000000000000,
24'b000000011011111111110011,
24'b111111111111000000000000,
24'b000000011100111111110010,
24'b000000000001000000000000,
24'b000000011101111111110100,
24'b000000000001000000000000,
24'b000000011101111111110100,
24'b000000000000111111111111,
24'b000000011110111111110100,
24'b000000000000000000000000,
24'b000000011111111111110100,
24'b111111111111000000000000,
24'b000000100000111111110011,
24'b111111111111000000000001,
24'b000000100000111111110011,
24'b111111111110000000000000,
24'b000000100000111111110001,
24'b000000000000111111111111,
24'b000000100010111111110001,
24'b000000000001000000000000,
24'b000000100011111111110001,
24'b000000000001111111111111,
24'b000000100101111111110010,
24'b000000000001000000000000,
24'b000000100110111111110010,
24'b000000000010000000000010,
24'b000000100101111111110100,
24'b111111111111000000000001,
24'b000000100110111111110000,
24'b000000000001000000000000,
24'b000000101001111111110010,
24'b000000000001000000000001,
24'b000000101001111111110010,
24'b000000000000000000000001,
24'b000000101010111111110010,
24'b111111111111000000000000,
24'b000000101101111111110001,
24'b000000000000000000000000,
24'b000000101111111111110001,
24'b111111111111000000000001,
24'b000000101111111111110000,
24'b000000000000000000000000,
24'b000000110010111111110000,
24'b111111111111000000000000,
24'b000000110100111111101110,
24'b000000000001000000000000,
24'b000000110111111111101111,
24'b000000000000000000000000,
24'b000000111010111111101111,
24'b000000000000000000000000,
24'b000000111101111111101110,
24'b000000000000000000000010,
24'b000000111111111111101101,
24'b000000000001000000000001,
24'b000001000010111111101110,
24'b111111111111000000000001,
24'b000001000100111111101011,
24'b000000000000111111111111,
24'b000001001011111111101011,
24'b111111111111000000000001,
24'b000001001110111111101000,
24'b000000000000000000000000,
24'b000001010100111111100111,
24'b111111111111000000000000,
24'b000001011001111111100100,
24'b000000000000111111111110,
24'b000001100010111111100000,
24'b000000000000111111111111,
24'b000001101010111111011100,
24'b000000000000111111111110,
24'b000001110110111111010101,
24'b000000000000000000000010,
24'b000001111101111111001011,
24'b000000000000000000000001,
24'b000010001001111110111010,
24'b000000000001111111111111,
24'b000010010110111110011100,
24'b111111111111000000000000,
24'b000010010011111101001111,
24'b000000000000000000000000,
24'b111111010001110111110100,
24'b001011010111110100101011,
24'b010100000100000010010001,
24'b001011010101001011010101,
24'b000110110011010000000111,
24'b110100101011001011010101,
24'b000001000001110111111110,
24'b001011010100001011010101,
24'b110100111111001110001010,
24'b110100101010110100101100,
24'b001111111001110111011010,
24'b001011010101001011010101,
24'b000100100010001110010010,
24'b110100101011001011010110,
24'b000000110001111000010000,
24'b001011010101001011010110,
24'b111101110000010000100000,
24'b110100101011001011010110,
24'b111001111011000010100001,
24'b110100101010001011010101,
24'b101110010111110100111010,
24'b001011010101110100101010,
24'b001000111011001111000000,
24'b110100101011001011010111,
24'b111011101110000010110100,
24'b110100101011001011010110,
24'b101110001101111101111101,
24'b110100101100110100101011,
24'b000111100110111000101100,
24'b110100101100001011010100,
24'b111001001011101010101100,
24'b001011010110001011010101,
24'b101001001100111010100011,
24'b001011010101110100101011,
24'b110111100110000010101110,
24'b001011010101110100101001,
24'b111101100000010010100010,
24'b110100101001110100101010,
24'b000011010010000100011010,
24'b110100101011110100101011,
24'b010001010110111111000010,
24'b110100101011001011010101,
24'b000000100110111001111110,
24'b110100101011001011010110,
24'b110000001100101101011111,
24'b001011010110110100101010,
24'b111111111100000111000101,
24'b110100101100110100101011,
24'b001111001001111000100111,
24'b110100101100001011010101,
24'b111000001001101000100010,
24'b001011010011110100101011,
24'b010000011000110110101101,
24'b001011010101001011010110,
24'b000011011001111100010011,
24'b001011010100001011010100,
24'b111110000110000001100011,
24'b001011010101001011010100,
24'b111000100001001110010111,
24'b110100101011001011010101,
24'b101010001101110101101110,
24'b001011010101110100101100,
24'b111001101100001011100100,
24'b110100101100110100101011,
24'b000001011001110100100000,
24'b001011010100110100101100,
24'b010000011000001010111001,
24'b110100101010001011010110,
24'b000000011010110100001000,
24'b001011010101001011010110,
24'b110001011100001010110101,
24'b110100101010110100101011,
24'b001001010010110100011101,
24'b001011010101001011010100,
24'b110011001010001100001111,
24'b110100101001110100101010,
24'b001010010010111101011100,
24'b110100101011001011010101,
24'b110100010010101110100101,
24'b001011010101110100101010,
24'b001100100101000101110111,
24'b110100101100001011010110,
24'b111110111110101110000111,
24'b001011010110001011010110,
24'b110111110011111100011100,
24'b001011010101001011010101,
24'b101000100101001010011001,
24'b110100101010110100101010,
24'b110111000100110000111011,
24'b001011010101110100101001,
24'b111100110101111110101111,
24'b001011010101110100101100,
24'b000010010011001100101111,
24'b110100101011110100101010,
24'b010000000010110100010001,
24'b001011010101001011010110,
24'b111110101110001001110001,
24'b110100101010001011010110,
24'b101101011100110001011101,
24'b001011010100110100101010,
24'b111011010110111111111101,
24'b001011010101110100101011,
24'b000001100110001111010010,
24'b110100101100110100101011,
24'b001110010101111110111100,
24'b110100101010001011010101,
24'b110100101010101111001101,
24'b001011010101110100101011,
24'b000010110000000101110100,
24'b110100101001110100101100,
24'b010001111111101101000101,
24'b001011010101001011010100,
24'b000001110001111001100011,
24'b001011010100001011010101,
24'b110010011000111110001000,
24'b001011010101110100101010,
24'b001001100010000010100010,
24'b001011010101001011010110,
24'b110001111000001110010011,
24'b110100101011110100101011,
24'b000000101111110011101010,
24'b001011010100110100101100,
24'b010000001100111111111011,
24'b001011010110001011010100,
24'b111111110000000110001000,
24'b001011010101001011010101,
24'b101111000101010100010101,
24'b110100101100110100101011,
24'b111101100111000100100011,
24'b110100101011110100101010,
24'b000100111101111100010110,
24'b110100101011110100101011,
24'b010100000011101100100001,
24'b001011010101001011010101,
24'b000101010010111010100110,
24'b001011010111001011010101,
24'b111111000011000000001010,
24'b001011010011001011010101,
24'b111000101101000101100011,
24'b001011010101001011010101,
24'b101001100100010011011000,
24'b110100101001110100101011,
24'b110111110011000010100000,
24'b110100101011110100101010,
24'b111100111100110010110000,
24'b001011010100110100101010,
24'b000000110110001001100010,
24'b110100101011110100101011,
24'b000101011000110001011111,
24'b001011010101110100101011,
24'b010001101100111111101010,
24'b001011010110001011010011,
24'b111000101001001101100101,
24'b110100101010110100101010,
24'b001101110101110100001100,
24'b001011010100001011010101,
24'b110101001001000010010010,
24'b001011010110110100101001,
24'b000010100110010001011010,
24'b110100101100110100101100,
24'b001001101100000000101110,
24'b110100101010110100101011,
24'b011001000100110000000000,
24'b001011010101001011010101,
24'b001010111111111111000110,
24'b001011010100001011010101,
24'b000110000101001101001101,
24'b110100101011001011010101,
24'b000010101001110011110100,
24'b001011010101001011010101,
24'b111111011000000001100110,
24'b001011010101001011010110,
24'b111010111101001111011100,
24'b110100101100001011010110,
24'b101101111001110110010001,
24'b001011010101110100101010,
24'b111111101111000100110011,
24'b001011010101110100101010,
24'b010001100011010100101111,
24'b110100101010001011010100,
24'b000100100001000110000010,
24'b110100101010001011010101,
24'b000000000111111111001001,
24'b110100101010001011010101,
24'b111100110101110001111000,
24'b001011010101001011010100,
24'b111001011110001011000100,
24'b110100101010001011010101,
24'b110100101010111100011001,
24'b110100101010001011010110,
24'b100110110100101100010101,
24'b001011010101110100101011,
24'b110111001000111010111110,
24'b001011010101110100101010,
24'b000101101111000010000001,
24'b001011010110001011010101,
24'b101100001101010000010101,
24'b110100101010110100101011,
24'b111000110011111111011001,
24'b110100101011110100101100,
24'b111110011001101110100100,
24'b001011010110110100101011,
24'b001010011101111101100001,
24'b001011010101001011010110,
24'b101111100110001011011000,
24'b110100101010110100101011,
24'b111011000101110001011110,
24'b001011010110110100101010,
24'b111111000010111101111110,
24'b001011010101110100101100,
24'b000010001101000011110101,
24'b001011010110110100101001,
24'b000110011001010000100111,
24'b110100101001110100101001,
24'b010010100100110111110000,
24'b001011010101001011010100,
24'b111001100000001101010110,
24'b110100101010110100101011,
24'b001111000100110101111001,
24'b001011010101001011010101,
24'b110111110010001011111000,
24'b110100101011110100101010,
24'b001110001001110100011100,
24'b001011010100001011010101,
24'b110111100000001001111101,
24'b110100101011110100101011,
24'b001110111101110001000001,
24'b001011010101001011010101,
24'b111111101011111101100001,
24'b001011010100001011010110,
24'b101111011001000010011100,
24'b001011010100110100101010,
24'b111110000110000111100011,
24'b001011010111110100101011,
24'b000101011011010101001101,
24'b110100101100110100101011,
24'b010100011010000100001000,
24'b110100101011001011010101,
24'b000101010000110011100001,
24'b001011010101001011010100,
24'b111101110001000011010000,
24'b001011010101001011010110,
24'b101110110111010011010101,
24'b110100101011110100101011,
24'b111110110111000100010010,
24'b110100101010110100101011,
24'b001101101010111100011100,
24'b110100101100001011010101,
24'b110101000000101100110000,
24'b001011010111110100101101,
24'b000011110101111010110010,
24'b001011010111110100101010,
24'b010100000010111111111000,
24'b001011010101001011010101,
24'b000101011110000011110101,
24'b001011010100001011010101,
24'b111110101010001000101011,
24'b001011010110001011010101,
24'b110001010000010110001011,
24'b110100101011110100101011,
24'b001001100100000100111000,
24'b110100101100001011010100,
24'b110011100100110011111000,
24'b001011010100110100101011,
24'b001010100000000010001011,
24'b001011010110001011010101,
24'b110011111100001001011001,
24'b001011010101110100101011,
24'b001010100110011000010010,
24'b110100101010001011010100,
24'b110011110101001000100110,
24'b110100101011110100101011,
24'b001010000101111010011111,
24'b001011010110001011010100,
24'b110010010010010100100010,
24'b110100101010110100101100,
24'b000001000110001000101011,
24'b110100101011110100101010,
24'b010000101100000100101111,
24'b110100101010001011010110,
24'b000000011000000001110110,
24'b110100101010001011010110,
24'b110000000100111110111110,
24'b110100101011110100101011,
24'b111111101010111011000100,
24'b110100101010110100101100,
24'b001110100101101111010000,
24'b001011010110001011010101,
24'b110111000010001001011000,
24'b110100101100110100101010,
24'b001110010010111011011001,
24'b110100101010001011010111,
24'b111110111100101011110110,
24'b001011010101001011010101,
24'b101110110110111010111001,
24'b001011010110110100101100,
24'b111110001110000010001110,
24'b001011010110110100101010,
24'b001100100100010000010000,
24'b110100101011001011010100,
24'b110011010011111000110101,
24'b001011010110110100101010,
24'b000001001010010000110111,
24'b110100101010110100101100,
24'b001110111101000011100100,
24'b110100101011001011010101,
24'b110101100110111101010101,
24'b110100101100110100101010,
24'b000011101011110000100010,
24'b001011010011110100101011,
24'b010010001010001001111111,
24'b110100101011001011010011,
24'b111010101011111011100111,
24'b110100101100110100101010,
24'b010010011011101011111000,
24'b001011010100001011010101,
24'b000100101101111010110101,
24'b001011010101001011010101,
24'b111101101111000010011000,
24'b001011010110001011010100,
24'b101111000111010001100000,
24'b110100101010110100101100,
24'b111111001101000010011100,
24'b110100101100110100101011,
24'b001110000100111011001011,
24'b110100101010001011010101,
24'b110101010111101101000100,
24'b001011010100110100101100,
24'b000100000100000100010000,
24'b110100101011110100101010,
24'b010011110001101011110100,
24'b001011010110001011010101,
24'b000011101111111000010001,
24'b001011010101001011010100,
24'b110011111111111100100100,
24'b001011010101110100101010,
24'b000100100001111111110100,
24'b001011010100110100101011,
24'b010101100001000011101010,
24'b001011010101001011010100,
24'b000111110100001111000011,
24'b110100101010001011010101,
24'b000010011111110011111011,
24'b001011010011001011010100,
24'b111101001110111111011010,
24'b001011010110001011010101,
24'b101111101001000011101101,
24'b001011010110110100101101,
24'b000000111000001000001110,
24'b001011010100110100101011,
24'b010001111000010100100001,
24'b110100101010001011010110,
24'b000010111010111011100011,
24'b001011010110001011010110,
24'b110100101101010001001111,
24'b110100101010110100101100,
24'b001101010101111010000010,
24'b001011010101001011010110,
24'b111000010000010000011110,
24'b110100101011110100101010,
24'b010001011101111001110100,
24'b001011010100001011010101,
24'b000101000010010000101101,
24'b110100101011001011010100,
24'b111111101001111010101110,
24'b001011010110001011010110,
24'b110011110011010011010000,
24'b110100101011110100101100,
24'b001110110100000110001011,
24'b110100101100001011010110,
24'b000011011100000000000010,
24'b110100101010001011010110,
24'b111111100101110011000101,
24'b001011010100001011010101,
24'b111100010101001011111011,
24'b110100101010001011010101,
24'b110111111011110110101000,
24'b001011010101001011010101,
24'b101010101100001111001101,
24'b110100101011110100101011,
24'b111011111100000001001111,
24'b110100101100110100101011,
24'b001100000100110011011101,
24'b001011010100001011010101,
24'b110101100110001100111000,
24'b110100101010110100101011,
24'b001110001011111110111011,
24'b110100101100001011010101,
24'b000001001111110000101011,
24'b001011010101001011010101,
24'b111011001011001000101000,
24'b110100101100001011010101,
24'b101110010000110010001110,
24'b001011010100110100101010,
24'b000110111110001000011000,
24'b110100101101001011010110,
24'b110001001101110000000000,
24'b001011010101110100101011,
24'b001000011000111100111000,
24'b001011010110001011010101,
24'b110010000000000010001010,
24'b001011010110110100101011,
24'b001000101101000111100000,
24'b001011010110001011010110,
24'b110001010101010100101111,
24'b110100101011110100101101,
24'b000000101100111101000100,
24'b001011010110110100101011,
24'b010001001010010101001011,
24'b110100101011001011010110,
24'b000010110000001000011100,
24'b110100101100001011010100,
24'b111011111010000011111101,
24'b110100101011001011010100,
24'b101101110010000000100011,
24'b110100101010110100101010,
24'b111110111011111101000000,
24'b110100101101110100101101,
24'b010000001001111000000111,
24'b110100101001001011010110,
24'b000010011111101001111110,
24'b001011010110001011010111,
24'b111101000100111001011010,
24'b001011010101001011010110,
24'b110111100100000000100110,
24'b001011010101001011010100,
24'b101001100111001101111111,
24'b110100101011110100101011,
24'b111010001010110100110101,
24'b001011010101110100101011,
24'b001001011110000011011001,
24'b001011010110001011010101,
24'b110001111000010011001001,
24'b110100101010110100101011,
24'b001000001010000011011100,
24'b110100101011001011010110,
24'b110001001001110100111011,
24'b001011010110110100101010,
24'b000111001111001101111110,
24'b110100101010001011010110,
24'b101111000110111111110000,
24'b110100101010110100101010,
24'b111101011000110001001111,
24'b001011010101110100101100,
24'b001011011010001000110110,
24'b110100101011001011010110,
24'b110010001111110001011100,
24'b001011010101110100101010,
24'b000000100111000000001001,
24'b001011010111110100101011,
24'b010000000001001110101001,
24'b110100101100001011010101,
24'b111111110111110101111100,
24'b001011010110001011010110,
24'b110000011011000100111100,
24'b001011010101110100101011,
24'b000111011100010101011001,
24'b110100101100001011010101,
24'b101111011001000111100000,
24'b110100101011110100101011,
24'b111100111000000010010101,
24'b110100101011110100101100,
24'b000011101100111110000101,
24'b110100101100110100101010,
24'b010010010000111000110000,
24'b110100101100001011010111,
24'b000001111110101010011000,
24'b001011010110001011010101,
24'b110010111010111001011010,
24'b001011010110110100101011,
24'b001010110010111111101000,
24'b001011010100001011010110,
24'b110100111101000101101010,
24'b001011010101110100101100,
24'b001101010010010100000101,
24'b110100101010001011010100,
24'b111111110010000011111000,
24'b110100101100001011010101,
24'b111000101101110100111011,
24'b001011010101001011010101,
24'b101001101011001100111100,
24'b110100101011110100101100,
24'b111000100001110111010000,
24'b001011010110110100101011,
24'b111111011000001111101001,
24'b110100101011110100101010,
24'b001100101100000001101010,
24'b110100101010001011010100,
24'b110100000111110011111100,
24'b001011010101110100101100,
24'b001001100010001101110000,
24'b110100101011001011010101,
24'b110001001011000000111101,
24'b110100101100110100101011,
24'b111111011010111010100100,
24'b110100101011110100101100,
24'b001101101111101100011001,
24'b001011010101001011010011,
24'b110101110111111101000101,
24'b001011010101110100101010,
24'b001100110100001101010100,
24'b110100101001001011010100,
24'b111101001100111101001000,
24'b110100101010001011010101,
24'b101100100100101100011111,
24'b001011010111110100101001,
24'b111010110011111010110010,
24'b001011010111110100101100,
24'b000001010011000001011000,
24'b001011010110110100101011,
24'b001110011011001110011101,
24'b110100101101001011010110,
24'b110101110001110101101010,
24'b001011010101110100101011,
24'b001011011010001010110001,
24'b110100101011001011010101,
24'b110011111100110001101111,
24'b001011010101110100101011,
24'b001001100110111110001111,
24'b001011010101001011010110,
24'b110000111111000011001011,
24'b001011010110110100101011,
24'b111110001011001000010011,
24'b001011010110110100101101,
24'b000100110011010101010000,
24'b110100101011110100101010,
24'b010011011000111101001100,
24'b001011010110001011010101,
24'b000011110100010100101001,
24'b110100101011001011010111,
24'b111011110010000110010000,
24'b110100101100001011010110,
24'b101100001011111000100001,
24'b001011010101110100101011,
24'b111010100110010010100101,
24'b110100101011110100101010,
24'b000001000001000110100101,
24'b110100101101110100101100,
24'b001101100111000010010001,
24'b110100101100001011010100,
24'b110011011110111110100100,
24'b110100101011110100101010,
24'b000000000110111001100110,
24'b110100101011110100101010,
24'b000110011110101011101000,
24'b001011010101110100101011,
24'b010100101101111011001110,
24'b001011010101001011010110,
24'b000100010011000010110001,
24'b001011010100001011010101,
24'b110101001111010000101101,
24'b110100101011110100101010,
24'b001101110001111000111101,
24'b001011010101001011010101,
24'b111110111000001111101000,
24'b110100101010001011010101,
24'b101110111100111001100110,
24'b001011010100110100101100,
24'b111110011100010001111011,
24'b110100101011110100101011,
24'b001100110101000100000010,
24'b110100101100001011010100,
24'b110011101010110110100010,
24'b001011010110110100101010,
24'b000001101001010000100001,
24'b110100101011110100101011,
24'b001111101010000011011011,
24'b110100101011001011010101,
24'b110110101000110110100110,
24'b001011010101110100101011,
24'b000101010111010001011110,
24'b110100101100110100101011,
24'b010101100100000110010100,
24'b110100101011001011010110,
24'b000111010101000011000001,
24'b110100101011001011010110,
24'b000001100110000000111000,
24'b110100101010001011010101,
24'b111011111101111111000100,
24'b110100101011001011010101,
24'b101110000000111101010011,
24'b110100101100110100101010,
24'b111110111001111011011011,
24'b110100101010110100101010,
24'b001111011010111001000000,
24'b110100101011001011010101,
24'b111111110100110101001110,
24'b110100101011001011010100,
24'b110000110000101001001001,
24'b001011010101110100101001,
24'b000111111111000001111000,
24'b110100101100001011010110,
24'b101111111110101011001000,
24'b001011010101110100101011,
24'b111101011100111010001111,
24'b001011010110110100101010,
24'b000011111111001001000010,
24'b110100101011110100101011,
24'b010001011010110001000011,
24'b001011010100001011010101,
24'b111001010010000110101111,
24'b110100101011110100101010,
24'b001111110011101110010001,
24'b001011010100001011010110,
24'b111001110001111011100000,
24'b001011010110110100101011,
24'b010010011111000010001011,
24'b001011010110001011010101,
24'b000110000011010000011010,
24'b110100101010001011010101,
24'b000001101001111111100101,
24'b110100101011001011010101,
24'b111110001111101111000000,
24'b001011010100001011010100,
24'b111010101100111110010111,
24'b001011010101001011010110,
24'b110101100110001101000000,
24'b110100101101001011010110,
24'b100111001111110100111110,
24'b001011010101110100101011,
24'b110110001010001010110011,
24'b110100101010110100101011,
24'b111100001001110010110000,
24'b001011010101110100101010,
24'b000001110100000001100000,
24'b001011010110110100101100,
24'b001111100100010001000111,
24'b110100101001001011010100,
24'b111110010011000000110100,
24'b110100101100001011010101,
24'b101100111101110000101001,
24'b001011010110110100101100,
24'b111010101000000000011101,
24'b001011010101110100101011,
24'b000000100101001111101010,
24'b110100101011110100101010,
24'b001100110001111000100100,
24'b001011010110001011010101,
24'b110010000000010000101001,
24'b110100101010110100101011,
24'b111101100100000011001101,
24'b110100101011110100101011,
24'b000001100001111100100011,
24'b110100101001110100101011,
24'b000100101011101110010010,
24'b001011010110110100101011,
24'b001000001001111111001011,
24'b001011010101110100101100,
24'b001101001111001111110001,
24'b110100101100110100101011,
24'b011011110000000000011000,
24'b110100101011001011010100,
24'b001101001111110001100111,
24'b001011010101001011010101,
24'b001000000101001001010011,
24'b110100101010001011010101,
24'b000100100011110010001011,
24'b001011010110001011010100,
24'b000001010101000001101011,
24'b001011010100001011010101,
24'b111101001101010001111011,
24'b110100101100001011010110,
24'b110001001100000010110000,
24'b110100101100110100101011,
24'b001010101010110100110011,
24'b001011010110001011010011,
24'b110110000001001110101101,
24'b110100101011110100101010,
24'b001111011100000010011011,
24'b110100101011001011010101,
24'b000011010011111101100000,
24'b110100101010001011010101,
24'b111110110011111000001010,
24'b110100101010001011010110,
24'b111010010011101010000101,
24'b001011010100001011010100,
24'b101110011000111001110011,
24'b001011010111110100101100,
24'b001000101110000001111010,
24'b001011010110001011010101,
24'b111011111110010001100100,
24'b110100101010001011010110,
24'b110101001010000011001101,
24'b110100101010001011010110,
24'b100101111100111101011000,
24'b110100101011110100101100,
24'b110100000101110111100010,
24'b110100101011110100101010,
24'b111001000000101001001001,
24'b001011010110110100101010,
24'b111100010100111001001001,
24'b001011010100110100101011,
24'b111111010101000111011100,
24'b110100101100110100101011,
24'b000011001000101101101010,
24'b001011010110110100101100,
24'b001110011110111001110000,
24'b001011010101001011010100,
24'b110011011100111110000000,
24'b001011010110110100101010,
24'b111111000010000001010101,
24'b001011010110110100101010,
24'b000011011011000100110111,
24'b001011010101110100101011,
24'b001000000110001001110111,
24'b001011010101110100101011,
24'b010100101011011000000011,
24'b110100101011001011010110,
24'b111100001101001000110011,
24'b110100101100110100101010,
24'b010011001110000001110011,
24'b110100101010001011010101,
24'b000100001101110100100001,
24'b001011010101001011010110,
24'b110101011000001101010101,
24'b110100101011110100101010,
24'b001101001100111000010111,
24'b001011010100001011010100,
24'b110110111010010001101010,
24'b110100101011110100101011,
24'b001101100101000101101011,
24'b110100101100001011010101,
24'b110110010001000001101011,
24'b110100101011110100101010,
24'b000101111000111110101101,
24'b110100101010110100101011,
24'b010110101111111011100111,
24'b110100101011001011010100,
24'b001001010010110111001111,
24'b110100101100001011010100,
24'b000100101101101010000100,
24'b001011010101001011010110,
24'b000001011001111011011100,
24'b001011010100001011010110,
24'b111110001001001100010011,
24'b110100101011001011010101,
24'b111001101011111100111010,
24'b110100101100001011010101,
24'b101100011101101101011111,
24'b001011010101110100101100,
24'b111101110111111110001001,
24'b001011010101110100101011,
24'b001110111001001111000111,
24'b110100101011001011010110,
24'b111111111001000001010000,
24'b110100101011001011010101,
24'b110001101110111011101000,
24'b110100101011110100101011,
24'b001010111000110101110101,
24'b110100101010001011010101,
24'b111100011111100111010001,
24'b001011010110001011010101,
24'b101101000001110110011111,
24'b001011010011110100101011,
24'b111101000100111101101110,
24'b001011010110110100101100,
24'b001100001101001100000101,
24'b110100101100001011010101,
24'b110100110001111011000000,
24'b110100101011110100101101,
24'b001011111011101001101000,
24'b001011010101001011010100,
24'b111100011011110110111100,
24'b001011010100001011010100,
24'b101011101110111011100110,
24'b001011010101110100101100,
24'b111001011100111111010000,
24'b001011010110110100101011,
24'b111110011011000011110111,
24'b001011010101110100101011,
24'b000010010101010000111110,
24'b110100101010110100101010,
24'b000111000010111111001111,
24'b110100101011110100101011,
24'b010011101101101101100010,
24'b001011010110001011010110,
24'b111011001111111010110101,
24'b001011010101110100101100,
24'b010001101101111111111111,
24'b001011010100001011010101,
24'b111110100100000111110000,
24'b111111111111000000000001,
24'b111111001110111100010000,
24'b001011010110110100101011,
24'b010100011100000101001001,
24'b001011010101001011010100,
24'b000111010010010010001111,
24'b110100101100001011010111,
24'b000001011110111001101001,
24'b001011010110001011010110,
24'b110101011010001111100010,
24'b110100101011110100101011,
24'b010000010011111000100100,
24'b001011010100001011010101,
24'b000100111001001111010000,
24'b110100101100001011010101,
24'b000001000111111001000110,
24'b001011010101001011010110,
24'b111110000100010001001111,
24'b110100101010001011010101,
24'b111010001110000011001000,
24'b110100101011001011010100,
24'b101110101010110101100000,
24'b001011010101110100101100,
24'b001001001001001111100001,
24'b110100101011001011010101,
24'b111011111101000011010010,
24'b110100101001001011010101,
24'b101110011100111110010110,
24'b110100101011110100101011,
24'b000111110101111001000011,
24'b110100101011001011010111,
24'b111001010101101011000001,
24'b001011010100001011010101,
24'b101001010110111010110101,
24'b001011010011110100101010,
24'b110111110010000010111101,
24'b001011010100110100101010,
24'b111101101010010010101110,
24'b110100101011110100101100,
24'b000011011001000100101001,
24'b110100101010110100101011,
24'b010001011111111111001101,
24'b110100101011001011010110,
24'b000000101101111010001010,
24'b110100101011001011010110,
24'b110000010100101101101001,
24'b001011010101110100101100,
24'b000000000001000111001110,
24'b110100101011110100101011,
24'b001111001111111000101110,
24'b110100101011001011010101,
24'b111000001110101000100110,
24'b001011010110110100101011,
24'b010000011110110110110100,
24'b001011010110001011010101,
24'b000011100000111100011010,
24'b001011010100001011010110,
24'b111110001011000001101000,
24'b001011010110001011010101,
24'b111000100101001110011101,
24'b110100101011001011010110,
24'b101010010000110101110010,
24'b001011010101110100101100,
24'b111001101110001011100111,
24'b110100101100110100101010,
24'b000001011100110100100010,
24'b001011010101110100101010,
24'b010000011100001010111100,
24'b110100101011001011010110,
24'b000000011101110100001011,
24'b001011010110001011010100,
24'b110001100000001010110111,
24'b110100101100110100101010,
24'b001001010110110100011111,
24'b001011011000001011010100,
24'b110011001101001100010011,
24'b110100101011110100101010,
24'b001010010100111101100010,
24'b110100101010001011010100,
24'b110100010111101110100111,
24'b001011010101110100101100,
24'b001100100101000101111010,
24'b110100101011001011010100,
24'b111111000010101110001001,
24'b001011010101001011010101,
24'b110111110111111100011110,
24'b001011010100001011010110,
24'b101000101000001010011001,
24'b110100101010110100101011,
24'b110111000110110000111011,
24'b001011010110110100101010,
24'b111100110101111110110000,
24'b001011010101110100101011,
24'b000010010100001100101111,
24'b110100101011110100101010,
24'b010000000010110100010001,
24'b001011010101001011010100,
24'b111110110000001001110001,
24'b110100101011001011010101,
24'b101101011111110001011110,
24'b001011010100110100101010,
24'b111011011000111111111100,
24'b001011010110110100101100,
24'b000001100111001111010011,
24'b110100101011110100101010,
24'b001110010111111110111011,
24'b110100101011001011010101,
24'b110100101011101111001101,
24'b001011010101110100101011,
24'b000010110001000101110010,
24'b110100101100110100101011,
24'b010010000001101101000110,
24'b001011010110001011010110,
24'b000001110001111001100011,
24'b001011010101001011010100,
24'b110010011001111110000111,
24'b001011010110110100101011,
24'b001001100010000010100011,
24'b001011010110001011010100,
24'b110001111010001110010101,
24'b110100101011110100101010,
24'b000000110001110011101010,
24'b001011010100110100101100,
24'b010000001110111111111100,
24'b001011010101001011010101,
24'b111111110000000110000111,
24'b001011010101001011010101,
24'b101111000101010100010110,
24'b110100101010110100101010,
24'b111101101000000100100010,
24'b110100101010110100101011,
24'b000100111100111100010110,
24'b110100101001110100101010,
24'b010100000011101100011111,
24'b001011010101001011010100,
24'b000101010011111010100101,
24'b001011010101001011010101,
24'b111111000100000000000110,
24'b001011010101001011010101,
24'b111000101101000101100010,
24'b001011010101001011010101,
24'b101001100100010011010110,
24'b110100101001110100101010,
24'b110111110101000010011111,
24'b110100101100110100101010,
24'b111100111110110010101111,
24'b001011010101110100101011,
24'b000000110110001001100011,
24'b110100101011110100101100,
24'b000101010111110001011111,
24'b001011010100110100101010,
24'b010001101110111111101000,
24'b001011010101001011010101,
24'b111000101001001101100001,
24'b110100101100110100101010,
24'b001101110110110100001011,
24'b001011010101001011010110,
24'b110101001010000010010010,
24'b001011010110110100101011,
24'b000010100100010001011010,
24'b110100101010110100101100,
24'b001001101101000000101100,
24'b110100101011110100101100,
24'b011001000011101111111111,
24'b001011010110001011010101,
24'b001010111110111111000110,
24'b001011010101001011010101,
24'b000110000011001101001101,
24'b110100101011001011010101,
24'b000010101001110011110100,
24'b001011010101001011010101,
24'b111111010111000001100110,
24'b001011010100001011010101,
24'b111010111100001111011011,
24'b110100101011001011010100,
24'b101101111100110110010000,
24'b001011010101110100101100,
24'b111111101110000100110001,
24'b001011010101110100101011,
24'b010001100010010100101110,
24'b110100101001001011010100,
24'b000100100001000110000000,
24'b110100101001001011010101,
24'b000000000101111111000111,
24'b110100101100001011010100,
24'b111100110110110001111001,
24'b001011010011001011010101,
24'b111001011101001011000011,
24'b110100101010001011010101,
24'b110100101001111100011000,
24'b110100101011001011010110,
24'b100110110010101100010100,
24'b001011010100110100101011,
24'b110111000111111010111100,
24'b001011010101110100101010,
24'b000101101110000001111111,
24'b001011010110001011010100,
24'b101100001101010000010100,
24'b110100101010110100101011,
24'b111000110010111111011000,
24'b110100101011110100101100,
24'b111110011000101110100011,
24'b001011010100110100101010,
24'b001010011100111101011111,
24'b001011010100001011010101,
24'b101111100110001011010101,
24'b110100101100110100101100,
24'b111011000110110001011101,
24'b001011010110110100101011,
24'b111111000001111101111101,
24'b001011010110110100101101,
24'b000010001101000011110100,
24'b001011010101110100101100,
24'b000110010111010000100110,
24'b110100101010110100101010,
24'b010010100010110111101110,
24'b001011010110001011010100,
24'b111001011111001101010101,
24'b110100101011110100101011,
24'b001111000010110101111010,
24'b001011010100001011010101,
24'b110111110001001011110111,
24'b110100101011110100101011,
24'b001110000111110100011010,
24'b001011010110001011010100,
24'b110111011110001001111101,
24'b110100101010110100101011,
24'b001110111011110000111111,
24'b001011010101001011010100,
24'b111111101010111101011111,
24'b001011010111001011010110,
24'b101111010111000010011100,
24'b001011010101110100101011,
24'b111110000011000111100101,
24'b001011010110110100101010,
24'b000101011010010101001101,
24'b110100101011110100101100,
24'b010100011000000100000111,
24'b110100101010001011010101,
24'b000101010000110011100000,
24'b001011010101001011010101,
24'b111101101110000011010000,
24'b001011010100001011010100,
24'b101110110111010011010101,
24'b110100101010110100101011,
24'b111110110101000100010010,
24'b110100101010110100101010,
24'b001101101001111100011011,
24'b110100101011001011010111,
24'b110100111100101100110000,
24'b001011010100110100101001,
24'b000011110111111010101111,
24'b001011010110110100101100,
24'b010011111111111111110100,
24'b001011010110001011010101,
24'b000101011101000011110011,
24'b001011010111001011010101,
24'b111110101000001000101100,
24'b001011010110001011010110,
24'b110001001110010110001011,
24'b110100101011110100101011,
24'b001001100011000100111000,
24'b110100101100001011010100,
24'b110011100010110011110110,
24'b001011010101110100101011,
24'b001010011110000010001011,
24'b001011010110001011010101,
24'b110011111100001001011001,
24'b001011010110110100101101,
24'b001010100100011000010010,
24'b110100101011001011010110,
24'b110011110011001000100110,
24'b110100101010110100101101,
24'b001010000010111010011110,
24'b001011010110001011010101,
24'b110010001110010100100000,
24'b110100101011110100101010,
24'b000001000101001000101011,
24'b110100101010110100101011,
24'b010000101001000100101101,
24'b110100101011001011010110,
24'b000000010100000001110110,
24'b110100101011001011010110,
24'b110000000000111110111110,
24'b110100101011110100101010,
24'b111111101000111011000100,
24'b110100101100110100101011,
24'b001110100011101111010010,
24'b001011010101001011010100,
24'b110111000001001001011000,
24'b110100101011110100101011,
24'b001110001111111011011001,
24'b110100101010001011010110,
24'b111110111011101011110101,
24'b001011010110001011010101,
24'b101110110011111010111010,
24'b001011010110110100101011,
24'b111110001110000010001111,
24'b001011010110110100101011,
24'b001100100010010000010000,
24'b110100101011001011010101,
24'b110011010001111000110101,
24'b001011010101110100101010,
24'b000001001000010000110111,
24'b110100101001110100101011,
24'b001110111100000011100010,
24'b110100101100001011010110,
24'b110101100100111101010101,
24'b110100101100110100101010,
24'b000011101010110000011111,
24'b001011010110110100101011,
24'b010010001000001010000000,
24'b110100101100001011010100,
24'b111010101000111011101001,
24'b110100101011110100101100,
24'b010010010110101011111000,
24'b001011010100001011010100,
24'b000100101011111010110110,
24'b001011010101001011010110,
24'b111101101011000010011001,
24'b001011010101001011010100,
24'b101111000011010001100000,
24'b110100101010110100101011,
24'b111111001011000010011101,
24'b110100101011110100101100,
24'b001101111111111011001010,
24'b110100101001001011010011,
24'b110101010101101101000011,
24'b001011010101110100101011,
24'b000100000010000100010001,
24'b110100101011110100101010,
24'b010011101110101011110101,
24'b001011010101001011010011,
24'b000011101111111000010010,
24'b001011010100001011010101,
24'b110011111101111100100100,
24'b001011010100110100101010,
24'b000100100000111111110100,
24'b001011010100110100101100,
24'b010101011111000011101010,
24'b001011010101001011010110,
24'b000111110001001111000010,
24'b110100101010001011010110,
24'b000010011100110011111010,
24'b001011010110001011010110,
24'b111101001001111111011100,
24'b001011010110001011010101,
24'b101111100100000011101110,
24'b001011010100110100101011,
24'b000000110101001000001100,
24'b001011010101110100101010,
24'b010001110101010100100001,
24'b110100101100001011010101,
24'b000010110111111011100101,
24'b001011010101001011010101,
24'b110100101011010001001110,
24'b110100101101110100101011,
24'b001101010100111010000100,
24'b001011010110001011010111,
24'b111000001100010000100000,
24'b110100101010110100101011,
24'b010001011001111001110100,
24'b001011010101001011010101,
24'b000100111110010000101110,
24'b110100101011001011010011,
24'b111111100110111010110000,
24'b001011010101001011010101,
24'b110011101111010011001111,
24'b110100101100110100101010,
24'b001110110001000110001100,
24'b110100101011001011010100,
24'b000011011001000000000001,
24'b110100101011001011010101,
24'b111111100011110011000111,
24'b001011010101001011010101,
24'b111100010010001011111100,
24'b110100101010001011010100,
24'b110111111000110110101010,
24'b001011010100001011010101,
24'b101010101010001111001100,
24'b110100101011110100101010,
24'b111011111011000001001111,
24'b110100101100110100101100,
24'b001100000001110011011110,
24'b001011010100001011010110,
24'b110101100011001100111000,
24'b110100101100110100101011,
24'b001110001000111110111101,
24'b110100101011001011010110,
24'b000001001011110000101011,
24'b001011011000001011010101,
24'b111011001000001000101100,
24'b110100101011001011010111,
24'b101110001011110010001111,
24'b001011010110110100101010,
24'b000110111001001000011101,
24'b110100101011001011010101,
24'b110001001010110000000001,
24'b001011010100110100101100,
24'b001000010100111100111010,
24'b001011010110001011010100,
24'b110001111110000010001011,
24'b001011010101110100101100,
24'b001000101000000111100001,
24'b001011010101001011010101,
24'b110001001111010100110001,
24'b110100101011110100101011,
24'b000000101001111101000101,
24'b001011010110110100101010,
24'b010001000111010101001101,
24'b110100101010001011010100,
24'b000010101110001000011111,
24'b110100101010001011010100,
24'b111011110111000011111100,
24'b110100101011001011010100,
24'b101101110000000000100011,
24'b110100101011110100101100,
24'b111110110111111101000011,
24'b110100101010110100101100,
24'b010000000111111000000101,
24'b110100101011001011010111,
24'b000010011010101010000000,
24'b001011010110001011010101,
24'b111101000010111001011011,
24'b001011010100001011010110,
24'b110111100010000000100111,
24'b001011010110001011010111,
24'b101001100001001110000001,
24'b110100101011110100101010,
24'b111010000111110100110110,
24'b001011010110110100101100,
24'b001001011010000011011011,
24'b001011010101001011010101,
24'b110001110100010011001010,
24'b110100101010110100101100,
24'b001000000101000011011110,
24'b110100101010001011010100,
24'b110001000110110100111100,
24'b001011010110110100101011,
24'b000111001010001101111110,
24'b110100101100001011010101,
24'b101111000011111111110010,
24'b110100101011110100101011,
24'b111101010100110001010000,
24'b001011010110110100101100,
24'b001011010110001000111010,
24'b110100101001001011010101,
24'b110010001011110001011100,
24'b001011010110110100101010,
24'b000000100010000000001101,
24'b001011010101110100101001,
24'b001111111111001110101001,
24'b110100101100001011010110,
24'b111111110010110101111101,
24'b001011010111001011010101,
24'b110000011000000100111110,
24'b001011010110110100101011,
24'b000111011000010101011011,
24'b110100101100001011010101,
24'b101111010100000111100010,
24'b110100101011110100101011,
24'b111100110011000010010111,
24'b110100101011110100101010,
24'b000011101001111110001000,
24'b110100101100110100101010,
24'b010010001011111000110100,
24'b110100101010001011010101,
24'b000001111011101010011010,
24'b001011010100001011010101,
24'b110010110101111001011010,
24'b001011010110110100101001,
24'b001010110000111111101010,
24'b001011010101001011010110,
24'b110100111000000101101101,
24'b001011010101110100101001,
24'b001101010001010100000111,
24'b110100101010001011010101,
24'b111111101111000011111011,
24'b110100101011001011010110,
24'b111000101010110100111110,
24'b001011010100001011010111,
24'b101001100101001100111110,
24'b110100101011110100101011,
24'b111000011100110111010010,
24'b001011010100110100101011,
24'b111111010101001111101011,
24'b110100101010110100101100,
24'b001100100110000001101001,
24'b110100101100001011010101,
24'b110100000000110011111111,
24'b001011010100110100101011,
24'b001001011101001101110001,
24'b110100101100001011010100,
24'b110001000101000001000001,
24'b110100101011110100101010,
24'b111111010110111010100111,
24'b110100101010110100101011,
24'b001101101101101100011011,
24'b001011010100001011010101,
24'b110101110011111101000110,
24'b001011010101110100101100,
24'b001100101100001101010110,
24'b110100101010001011010011,
24'b111101000111111101001100,
24'b110100101010001011010101,
24'b101100011110101100100011,
24'b001011010101110100101010,
24'b111010101101111010110101,
24'b001011010101110100101100,
24'b000001001101000001011000,
24'b001011010111110100101010,
24'b001110010110001110100001,
24'b110100101010001011010110,
24'b110101101011110101101010,
24'b001011010110110100101011,
24'b001011010101001010110011,
24'b110100101100001011010101,
24'b110011110110110001110001,
24'b001011010101110100101010,
24'b001001100001111110010010,
24'b001011010101001011010101,
24'b110000111010000011001111,
24'b001011010101110100101100,
24'b111110000100001000010100,
24'b001011010110110100101010,
24'b000100110001010101010011,
24'b110100101011110100101101,
24'b010011010001111101001111,
24'b001011010110001011010101,
24'b000011101110010100101011,
24'b110100101011001011010110,
24'b111011101110000110010010,
24'b110100101100001011010110,
24'b101100000101111000100011,
24'b001011010111110100101010,
24'b111010100001010010101010,
24'b110100101100110100101011,
24'b000000111011000110101010,
24'b110100101010110100101100,
24'b001101100010000010010100,
24'b110100101010001011010101,
24'b110011011001111110100101,
24'b110100101011110100101100,
24'b111111111111111001101001,
24'b110100101011110100101010,
24'b000110010111101011101001,
24'b001011010110110100101011,
24'b010100100111111011010010,
24'b001011010101001011010101,
24'b000100001101000010110011,
24'b001011010101001011010100,
24'b110101001010010000110010,
24'b110100101010110100101011,
24'b001101101010111001000000,
24'b001011010110001011010101,
24'b111110110010001111101100,
24'b110100101010001011010110,
24'b101110110101111001101010,
24'b001011010011110100101100,
24'b111110010110010001111110,
24'b110100101011110100101100,
24'b001100101111000100000111,
24'b110100101011001011010101,
24'b110011100011110110100111,
24'b001011010101110100101011,
24'b000001100000010000100100,
24'b110100101011110100101010,
24'b001111100100000011011111,
24'b110100101100001011010110,
24'b110110100001110110101010,
24'b001011010101110100101100,
24'b000101001111010001100010,
24'b110100101011110100101011,
24'b010101011100000110010110,
24'b110100101100001011010110,
24'b000111001100000011000101,
24'b110100101010001011010100,
24'b000001100000000000111011,
24'b110100101011001011010110,
24'b111011110110111111001000,
24'b110100101011001011010110,
24'b101101111000111101011000,
24'b110100101010110100101010,
24'b111110110001111011011101,
24'b110100101100110100101011,
24'b001111010001111001000100,
24'b110100101011001011010101,
24'b111111101100110101010011,
24'b110100101010001011010101,
24'b110000100111101001001101,
24'b001011010101110100101010,
24'b000111110110000001111100,
24'b110100101101001011010110,
24'b101111110110101011001100,
24'b001011010110110100101001,
24'b111101010100111010010100,
24'b001011010101110100101001,
24'b000011111001001001000110,
24'b110100101011110100101101,
24'b010001010001110001000101,
24'b001011010110001011010110,
24'b111001001001000110110100,
24'b110100101011110100101010,
24'b001111101010101110010100,
24'b001011010110001011010110,
24'b111001101000111011100111,
24'b001011010110110100101011,
24'b010010010110000010010000,
24'b001011010110001011010101,
24'b000101111001010000011111,
24'b110100101100001011010101,
24'b000001100000111111101011,
24'b110100101010001011010110,
24'b111110000101101111000101,
24'b001011010100001011010100,
24'b111010100001111110011101,
24'b001011010101001011010101,
24'b110101011011001101001000,
24'b110100101011001011010100,
24'b100111000111110101000100,
24'b001011010100110100101100,
24'b110110000010001010110111,
24'b110100101011110100101101,
24'b111011111110110010110110,
24'b001011010101110100101011,
24'b000001101001000001101000,
24'b001011010011110100101010,
24'b001111011011010001001010,
24'b110100101010001011010101,
24'b111110000111000000111010,
24'b110100101010001011010101,
24'b101100110001110000101101,
24'b001011010111110100101011,
24'b111010011101000000100011,
24'b001011010101110100101010,
24'b000000011010001111110000,
24'b110100101011110100101010,
24'b001100100110111000101011,
24'b001011010011001011010110,
24'b110001110101010000101101,
24'b110100101010110100101011,
24'b111101011000000011010010,
24'b110100101100110100101001,
24'b000001010110111100101001,
24'b110100101001110100101010,
24'b000100011111101110011001,
24'b001011010101110100101010,
24'b000111111111111111010000,
24'b001011010100110100101011,
24'b001101000100001111110110,
24'b110100101011110100101011,
24'b011011100101000000011101,
24'b110100101011001011010101,
24'b001101000010110001101101,
24'b001011010100001011010110,
24'b000111111001001001011001,
24'b110100101011001011010101,
24'b000100010110110010010011,
24'b001011010100001011010101,
24'b000001000111000001101111,
24'b001011010101001011010100,
24'b111101000000010010000010,
24'b110100101011001011010110,
24'b110000111111000010111000,
24'b110100101001110100101011,
24'b001010011110110100110111,
24'b001011010101001011010110,
24'b110101110001001110110001,
24'b110100101100110100101011,
24'b001111001100000010100000,
24'b110100101100001011010101,
24'b000011000011111101100111,
24'b110100101010001011010101,
24'b111110100001111000001111,
24'b110100101100001011010100,
24'b111010000101101010001100,
24'b001011010110001011010110,
24'b101110001000111001111101,
24'b001011010101110100101100,
24'b001000011101000010000000,
24'b001011010110001011010110,
24'b111011101110010001101010,
24'b110100101100001011010110,
24'b110100111000000011010110,
24'b110100101010001011010110,
24'b100101101001111101011111,
24'b110100101100110100101010,
24'b110011110100110111101010,
24'b110100101100110100101001,
24'b111000101110101001010010,
24'b001011010101110100101011,
24'b111100000001111001010000,
24'b001011010110110100101010,
24'b111111000001000111100110,
24'b110100101011110100101010,
24'b000010110101101101110010,
24'b001011010110110100101010,
24'b001110001101111001111001,
24'b001011010110001011010110,
24'b110011000111111110001011,
24'b001011010011110100101100,
24'b111110101101000001011011,
24'b001011010110110100101100,
24'b000011000011000100111110,
24'b001011010110110100101010,
24'b000111101111001001111111,
24'b001011010110110100101100,
24'b010100010100011000001101,
24'b110100101010001011010110,
24'b111011110111001000111101,
24'b110100101001110100101011,
24'b010010110101000001111001,
24'b110100101100001011010111,
24'b000011110010110100101001,
24'b001011010111001011010101,
24'b110101000000001101100000,
24'b110100101011110100101011,
24'b001100110010111000100000,
24'b001011010101001011010110,
24'b110110011101010001110101,
24'b110100101010110100101010,
24'b001101001010000101110101,
24'b110100101011001011010111,
24'b110101110011000001110101,
24'b110100101011110100101011,
24'b000101011001111110110111,
24'b110100101010110100101011,
24'b010110010001111011110010,
24'b110100101011001011010110,
24'b001000110000110111011011,
24'b110100101010001011010110,
24'b000100000111101010001101,
24'b001011010100001011010101,
24'b000000110110111011100110,
24'b001011010101001011010110,
24'b111101100100001100100000,
24'b110100101001001011010110,
24'b111001000100111101000100,
24'b110100101100001011010101,
24'b101011110011101101101010,
24'b001011010101110100101001,
24'b111101001111111110010101,
24'b001011010100110100101010,
24'b001110001110001111010100,
24'b110100101010001011010101,
24'b111111001101000001011100,
24'b110100101010001011010101,
24'b110000111111111011110100,
24'b110100101001110100101011,
24'b001010000111110101111111,
24'b110100101011001011010110,
24'b111011101010100111011110,
24'b001011010111001011010101,
24'b101100001001110110101110,
24'b001011010101110100101010,
24'b111100001010111110000000,
24'b001011010101110100101100,
24'b001011010000001100010111,
24'b110100101000001011010101,
24'b110011101110111011001110,
24'b110100101011110100101001,
24'b001010111001101001111000,
24'b001011010101001011010101,
24'b111011010010110111001111,
24'b001011010101001011010101,
24'b101010011110111011111011,
24'b001011010110110100101011,
24'b111000000111111111101010,
24'b001011010101110100101010,
24'b111100111111000100010001,
24'b001011010110110100101011,
24'b000000110010010001011110,
24'b110100101011110100101011,
24'b000101010101111111110110,
24'b110100101010110100101011,
24'b010001110100101110010100,
24'b001011010100001011010101,
24'b111001001011111011110110,
24'b001011010100110100101011,
24'b001111011111000001100000,
24'b001011010100001011010110,
24'b111100010110001010011100,
24'b000000000000000000000001,
24'b000000000100000100011000,
24'b000000000000000000000000,
24'b000000100000000010110101,
24'b000000000000000000000001,
24'b000000100100000010000101,
24'b000000000001000000000000,
24'b000000100100000001101000,
24'b111111111111000000000000,
24'b000000100010000001010011,
24'b000000000001000000000000,
24'b000000011111000001000110,
24'b111111111111000000000000,
24'b000000011100000000111001,
24'b000000000000111111111110,
24'b000000011101000000110001,
24'b000000000001111111111111,
24'b000000011011000000101100,
24'b111111111111111111111111,
24'b000000011010000000100101,
24'b111111111111000000000000,
24'b000000011000000000100000,
24'b111111111111000000000001,
24'b000000010110000000011011,
24'b000000000000000000000000,
24'b000000010110000000010111,
24'b000000000001000000000001,
24'b000000010100000000010110,
24'b000000000000000000000001,
24'b000000010010000000010011,
24'b000000000000000000000001,
24'b000000010001000000010001,
24'b000000000000000000000000,
24'b000000010001000000001111,
24'b111111111111000000000001,
24'b000000001111000000001100,
24'b000000000001000000000000,
24'b000000001111000000001101,
24'b111111111111111111111111,
24'b000000001111000000001001,
24'b000000000000111111111111,
24'b000000001111000000001001,
24'b000000000000000000000000,
24'b000000001110000000000111,
24'b000000000000000000000000,
24'b000000001101000000000110,
24'b000000000000111111111111,
24'b000000001110000000000101,
24'b000000000001111111111111,
24'b000000001110000000000110,
24'b111111111111000000000000,
24'b000000001101000000000011,
24'b000000000000111111111111,
24'b000000001101000000000011,
24'b000000000000111111111111,
24'b000000001101000000000010,
24'b000000000001000000000000,
24'b000000001101000000000011,
24'b111111111110000000000000,
24'b000000001100000000000001,
24'b111111111111000000000000,
24'b000000001100000000000000,
24'b111111111111000000000000,
24'b000000001100000000000000,
24'b111111111111000000000000,
24'b000000001011111111111111,
24'b000000000000000000000000,
24'b000000001011111111111111,
24'b000000000001000000000000,
24'b000000001100000000000000,
24'b111111111111000000000001,
24'b000000001001111111111110,
24'b111111111111111111111111,
24'b000000001011111111111101,
24'b000000000001000000000000,
24'b000000001011111111111110,
24'b000000000000000000000000,
24'b000000001011111111111111,
24'b111111111111000000000000,
24'b000000001010111111111110,
24'b111111111110000000000000,
24'b000000001001111111111011,
24'b000000000000111111111111,
24'b000000001010111111111100,
24'b000000000001111111111111,
24'b000000001011111111111101,
24'b000000000000000000000000,
24'b000000001011111111111101,
24'b111111111110000000000000,
24'b000000001011111111111010,
24'b000000000001000000000000,
24'b000000001010111111111100,
24'b000000000000000000000000,
24'b000000001010111111111010,
24'b000000000010000000000000,
24'b000000001010111111111101,
24'b000000000001000000000001,
24'b000000001010111111111101,
24'b000000000000000000000001,
24'b000000001000111111111011,
24'b000000000001111111111111,
24'b000000001001111111111100,
24'b000000000000000000000000,
24'b000000001001111111111100,
24'b000000000000111111111110,
24'b000000001010111111111100,
24'b000000000000111111111111,
24'b000000001011111111111011,
24'b000000000000000000000000,
24'b000000001011111111111011,
24'b000000000001000000000001,
24'b000000001010111111111100,
24'b000000000000000000000001,
24'b000000001010111111111011,
24'b000000000000000000000001,
24'b000000001001111111111011,
24'b000000000000000000000001,
24'b000000001000111111111011,
24'b000000000000111111111111,
24'b000000001010111111111011,
24'b000000000000000000000001,
24'b000000000111111111111010,
24'b000000000001111111111111,
24'b000000001010111111111011,
24'b000000000001000000000000,
24'b000000001000111111111100,
24'b111111111111111111111111,
24'b000000001010111111111010,
24'b000000000000000000000001,
24'b000000001000111111111010,
24'b000000000000111111111110,
24'b000000001010111111111010,
24'b000000000000000000000000,
24'b000000001010111111111001,
24'b000000000010000000000001,
24'b000000001001111111111100,
24'b111111111111000000000000,
24'b000000001010111111111010,
24'b000000000000000000000000,
24'b000000001010111111111010,
24'b000000000000000000000010,
24'b000000001001111111111010,
24'b000000000001000000000001,
24'b000000001001111111111011,
24'b111111111111000000000000,
24'b000000001000111111111001,
24'b000000000001000000000000,
24'b000000001001111111111011,
24'b111111111111000000000000,
24'b000000001010111111111001,
24'b000000000001000000000001,
24'b000000001000111111111010,
24'b000000000000000000000000,
24'b000000001001111111111001,
24'b000000000001000000000000,
24'b000000001010111111111011,
24'b000000000000000000000001,
24'b000000001001111111111010,
24'b000000000000000000000001,
24'b000000000111111111111011,
24'b000000000000111111111111,
24'b000000001001111111111010,
24'b000000000000111111111111,
24'b000000001010111111111010,
24'b000000000000000000000001,
24'b000000001001111111111011,
24'b111111111111000000000001,
24'b000000001000111111111010,
24'b111111111111111111111111,
24'b000000001010111111111001,
24'b000000000000000000000001,
24'b000000001000111111111001,
24'b000000000000111111111111,
24'b000000001010111111111010,
24'b000000000000000000000001,
24'b000000001001111111111010,
24'b000000000000000000000000,
24'b000000001001111111111010,
24'b111111111111000000000000,
24'b000000001010111111111001,
24'b000000000000000000000001,
24'b000000001001111111111010,
24'b000000000000000000000001,
24'b000000001000111111111010,
24'b111111111111111111111111,
24'b000000001010111111111010,
24'b111111111111000000000000,
24'b000000001001111111111001,
24'b000000000001000000000000,
24'b000000001010111111111010,
24'b000000000000000000000001,
24'b000000001001111111111011,
24'b111111111110000000000000,
24'b000000001010111111111000,
24'b000000000000000000000000,
24'b000000001010111111111001,
24'b111111111111000000000001,
24'b000000001010111111111000,
24'b000000000001000000000001,
24'b000000001001111111111010,
24'b000000000001000000000001,
24'b000000001001111111111010,
24'b000000000001000000000001,
24'b000000001000111111111011,
24'b111111111111000000000000,
24'b000000001000111111111001,
24'b000000000000111111111111,
24'b000000001010111111111001,
24'b000000000001000000000000,
24'b000000001010111111111010,
24'b111111111111000000000010,
24'b000000001000111111111000,
24'b000000000000000000000000,
24'b000000001000111111111010,
24'b111111111110111111111111,
24'b000000001010111111110111,
24'b000000000001000000000000,
24'b000000001001111111111001,
24'b111111111111000000000000,
24'b000000001010111111111000,
24'b000000000000000000000000,
24'b000000001010111111111000,
24'b000000000010000000000001,
24'b000000001001111111111010,
24'b000000000000111111111111,
24'b000000001011111111111001,
24'b000000000001000000000001,
24'b000000001010111111111010,
24'b111111111111000000000001,
24'b000000001001111111111001,
24'b000000000000000000000000,
24'b000000001010111111111010,
24'b111111111111000000000001,
24'b000000001001111111111000,
24'b000000000000000000000001,
24'b000000001000111111111000,
24'b000000000000111111111110,
24'b000000001011111111111000,
24'b000000000001000000000000,
24'b000000001010111111111001,
24'b000000000000000000000000,
24'b000000001011111111111001};